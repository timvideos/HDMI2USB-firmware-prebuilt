/* Machine-generated using LiteX gen */
module top(
	input clk100,
	input cpu_reset,
	output reg serial_tx,
	input serial_rx,
	input user_sw0,
	output oled_dc,
	output oled_res,
	output oled_sclk,
	output oled_sdin,
	output oled_vbat,
	output oled_vdd,
	output [14:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output [1:0] ddram_dm,
	inout [15:0] ddram_dq,
	output [1:0] ddram_dqs_p,
	output [1:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output reg spiflash_1x_cs_n,
	output reg spiflash_1x_mosi,
	input spiflash_1x_miso,
	output spiflash_1x_wp,
	output spiflash_1x_hold,
	output eth_clocks_tx,
	input eth_clocks_rx,
	output eth_rst_n,
	input eth_int_n,
	inout eth_mdio,
	output eth_mdc,
	input eth_rx_ctl,
	input [3:0] eth_rx_data,
	output eth_tx_ctl,
	output [3:0] eth_tx_data,
	input hdmi_in_clk_p,
	input hdmi_in_clk_n,
	input hdmi_in_data0_p,
	input hdmi_in_data0_n,
	input hdmi_in_data1_p,
	input hdmi_in_data1_n,
	input hdmi_in_data2_p,
	input hdmi_in_data2_n,
	input hdmi_in_scl,
	inout hdmi_in_sda,
	output hdmi_in_hpd_en,
	input hdmi_in_cec,
	output hdmi_in_txen,
	output hdmi_out_clk_p,
	output hdmi_out_clk_n,
	output hdmi_out_data0_p,
	output hdmi_out_data0_n,
	output hdmi_out_data1_p,
	output hdmi_out_data1_n,
	output hdmi_out_data2_p,
	output hdmi_out_data2_n,
	input hdmi_out_scl,
	input hdmi_out_sda,
	input hdmi_out_cec,
	input hdmi_out_hdp
);

wire [29:0] videosoc_videosoc_ibus_adr;
wire [31:0] videosoc_videosoc_ibus_dat_w;
wire [31:0] videosoc_videosoc_ibus_dat_r;
wire [3:0] videosoc_videosoc_ibus_sel;
wire videosoc_videosoc_ibus_cyc;
wire videosoc_videosoc_ibus_stb;
wire videosoc_videosoc_ibus_ack;
wire videosoc_videosoc_ibus_we;
wire [2:0] videosoc_videosoc_ibus_cti;
wire [1:0] videosoc_videosoc_ibus_bte;
wire videosoc_videosoc_ibus_err;
wire [29:0] videosoc_videosoc_dbus_adr;
wire [31:0] videosoc_videosoc_dbus_dat_w;
wire [31:0] videosoc_videosoc_dbus_dat_r;
wire [3:0] videosoc_videosoc_dbus_sel;
wire videosoc_videosoc_dbus_cyc;
wire videosoc_videosoc_dbus_stb;
wire videosoc_videosoc_dbus_ack;
wire videosoc_videosoc_dbus_we;
wire [2:0] videosoc_videosoc_dbus_cti;
wire [1:0] videosoc_videosoc_dbus_bte;
wire videosoc_videosoc_dbus_err;
reg [31:0] videosoc_videosoc_interrupt = 32'd0;
wire [31:0] videosoc_videosoc_i_adr_o;
wire [31:0] videosoc_videosoc_d_adr_o;
wire [29:0] videosoc_videosoc_rom_bus_adr;
wire [31:0] videosoc_videosoc_rom_bus_dat_w;
wire [31:0] videosoc_videosoc_rom_bus_dat_r;
wire [3:0] videosoc_videosoc_rom_bus_sel;
wire videosoc_videosoc_rom_bus_cyc;
wire videosoc_videosoc_rom_bus_stb;
reg videosoc_videosoc_rom_bus_ack = 1'd0;
wire videosoc_videosoc_rom_bus_we;
wire [2:0] videosoc_videosoc_rom_bus_cti;
wire [1:0] videosoc_videosoc_rom_bus_bte;
reg videosoc_videosoc_rom_bus_err = 1'd0;
wire [12:0] videosoc_videosoc_rom_adr;
wire [31:0] videosoc_videosoc_rom_dat_r;
wire [29:0] videosoc_videosoc_sram_bus_adr;
wire [31:0] videosoc_videosoc_sram_bus_dat_w;
wire [31:0] videosoc_videosoc_sram_bus_dat_r;
wire [3:0] videosoc_videosoc_sram_bus_sel;
wire videosoc_videosoc_sram_bus_cyc;
wire videosoc_videosoc_sram_bus_stb;
reg videosoc_videosoc_sram_bus_ack = 1'd0;
wire videosoc_videosoc_sram_bus_we;
wire [2:0] videosoc_videosoc_sram_bus_cti;
wire [1:0] videosoc_videosoc_sram_bus_bte;
reg videosoc_videosoc_sram_bus_err = 1'd0;
wire [12:0] videosoc_videosoc_sram_adr;
wire [31:0] videosoc_videosoc_sram_dat_r;
reg [3:0] videosoc_videosoc_sram_we = 4'd0;
wire [31:0] videosoc_videosoc_sram_dat_w;
reg [13:0] videosoc_videosoc_interface_adr = 14'd0;
reg videosoc_videosoc_interface_we = 1'd0;
reg [7:0] videosoc_videosoc_interface_dat_w = 8'd0;
wire [7:0] videosoc_videosoc_interface_dat_r;
wire [29:0] videosoc_videosoc_bus_wishbone_adr;
wire [31:0] videosoc_videosoc_bus_wishbone_dat_w;
reg [31:0] videosoc_videosoc_bus_wishbone_dat_r = 32'd0;
wire [3:0] videosoc_videosoc_bus_wishbone_sel;
wire videosoc_videosoc_bus_wishbone_cyc;
wire videosoc_videosoc_bus_wishbone_stb;
reg videosoc_videosoc_bus_wishbone_ack = 1'd0;
wire videosoc_videosoc_bus_wishbone_we;
wire [2:0] videosoc_videosoc_bus_wishbone_cti;
wire [1:0] videosoc_videosoc_bus_wishbone_bte;
reg videosoc_videosoc_bus_wishbone_err = 1'd0;
reg [1:0] videosoc_videosoc_counter = 2'd0;
reg [31:0] videosoc_videosoc_load_storage_full = 32'd0;
wire [31:0] videosoc_videosoc_load_storage;
reg videosoc_videosoc_load_re = 1'd0;
reg [31:0] videosoc_videosoc_reload_storage_full = 32'd0;
wire [31:0] videosoc_videosoc_reload_storage;
reg videosoc_videosoc_reload_re = 1'd0;
reg videosoc_videosoc_en_storage_full = 1'd0;
wire videosoc_videosoc_en_storage;
reg videosoc_videosoc_en_re = 1'd0;
wire videosoc_videosoc_update_value_re;
wire videosoc_videosoc_update_value_r;
reg videosoc_videosoc_update_value_w = 1'd0;
reg [31:0] videosoc_videosoc_value_status = 32'd0;
wire videosoc_videosoc_irq;
wire videosoc_videosoc_zero_status;
reg videosoc_videosoc_zero_pending = 1'd0;
wire videosoc_videosoc_zero_trigger;
reg videosoc_videosoc_zero_clear = 1'd0;
reg videosoc_videosoc_zero_old_trigger = 1'd0;
wire videosoc_videosoc_eventmanager_status_re;
wire videosoc_videosoc_eventmanager_status_r;
wire videosoc_videosoc_eventmanager_status_w;
wire videosoc_videosoc_eventmanager_pending_re;
wire videosoc_videosoc_eventmanager_pending_r;
wire videosoc_videosoc_eventmanager_pending_w;
reg videosoc_videosoc_eventmanager_storage_full = 1'd0;
wire videosoc_videosoc_eventmanager_storage;
reg videosoc_videosoc_eventmanager_re = 1'd0;
reg [31:0] videosoc_videosoc_value = 32'd0;
wire [29:0] videosoc_interface0_wb_sdram_adr;
wire [31:0] videosoc_interface0_wb_sdram_dat_w;
reg [31:0] videosoc_interface0_wb_sdram_dat_r = 32'd0;
wire [3:0] videosoc_interface0_wb_sdram_sel;
wire videosoc_interface0_wb_sdram_cyc;
wire videosoc_interface0_wb_sdram_stb;
reg videosoc_interface0_wb_sdram_ack = 1'd0;
wire videosoc_interface0_wb_sdram_we;
wire [2:0] videosoc_interface0_wb_sdram_cti;
wire [1:0] videosoc_interface0_wb_sdram_bte;
reg videosoc_interface0_wb_sdram_err = 1'd0;
(* dont_touch = "true" *) wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire sys4x_dqs_clk;
wire clk200_clk;
wire clk200_rst;
wire clk100_clk;
wire clk100_rst;
wire videosoc_pll_locked;
wire videosoc_pll_fb;
wire videosoc_pll_sys;
wire videosoc_pll_sys4x;
wire videosoc_pll_sys4x_dqs;
wire videosoc_pll_clk200;
reg [3:0] videosoc_reset_counter = 4'd15;
reg videosoc_ic_reset = 1'd1;
wire videosoc_rs232phyinterface0_sink_valid;
reg videosoc_rs232phyinterface0_sink_ready = 1'd0;
wire videosoc_rs232phyinterface0_sink_first;
wire videosoc_rs232phyinterface0_sink_last;
wire [7:0] videosoc_rs232phyinterface0_sink_payload_data;
reg videosoc_rs232phyinterface0_source_valid = 1'd0;
wire videosoc_rs232phyinterface0_source_ready;
reg videosoc_rs232phyinterface0_source_first = 1'd0;
reg videosoc_rs232phyinterface0_source_last = 1'd0;
reg [7:0] videosoc_rs232phyinterface0_source_payload_data = 8'd0;
reg videosoc_rs232phyinterface1_sink_valid = 1'd0;
reg videosoc_rs232phyinterface1_sink_ready = 1'd0;
reg videosoc_rs232phyinterface1_sink_first = 1'd0;
wire videosoc_rs232phyinterface1_sink_last;
reg [7:0] videosoc_rs232phyinterface1_sink_payload_data = 8'd0;
reg videosoc_rs232phyinterface1_source_valid = 1'd0;
wire videosoc_rs232phyinterface1_source_ready;
reg videosoc_rs232phyinterface1_source_first = 1'd0;
reg videosoc_rs232phyinterface1_source_last = 1'd0;
reg [7:0] videosoc_rs232phyinterface1_source_payload_data = 8'd0;
wire videosoc_uart_rxtx_re;
wire [7:0] videosoc_uart_rxtx_r;
wire [7:0] videosoc_uart_rxtx_w;
wire videosoc_uart_txfull_status;
wire videosoc_uart_rxempty_status;
wire videosoc_uart_irq;
wire videosoc_uart_tx_status;
reg videosoc_uart_tx_pending = 1'd0;
wire videosoc_uart_tx_trigger;
reg videosoc_uart_tx_clear = 1'd0;
reg videosoc_uart_tx_old_trigger = 1'd0;
wire videosoc_uart_rx_status;
reg videosoc_uart_rx_pending = 1'd0;
wire videosoc_uart_rx_trigger;
reg videosoc_uart_rx_clear = 1'd0;
reg videosoc_uart_rx_old_trigger = 1'd0;
wire videosoc_uart_status_re;
wire [1:0] videosoc_uart_status_r;
reg [1:0] videosoc_uart_status_w = 2'd0;
wire videosoc_uart_pending_re;
wire [1:0] videosoc_uart_pending_r;
reg [1:0] videosoc_uart_pending_w = 2'd0;
reg [1:0] videosoc_uart_storage_full = 2'd0;
wire [1:0] videosoc_uart_storage;
reg videosoc_uart_re = 1'd0;
wire videosoc_uart_tx_fifo_sink_valid;
wire videosoc_uart_tx_fifo_sink_ready;
reg videosoc_uart_tx_fifo_sink_first = 1'd0;
reg videosoc_uart_tx_fifo_sink_last = 1'd0;
wire [7:0] videosoc_uart_tx_fifo_sink_payload_data;
wire videosoc_uart_tx_fifo_source_valid;
wire videosoc_uart_tx_fifo_source_ready;
wire videosoc_uart_tx_fifo_source_first;
wire videosoc_uart_tx_fifo_source_last;
wire [7:0] videosoc_uart_tx_fifo_source_payload_data;
wire videosoc_uart_tx_fifo_syncfifo_we;
wire videosoc_uart_tx_fifo_syncfifo_writable;
wire videosoc_uart_tx_fifo_syncfifo_re;
wire videosoc_uart_tx_fifo_syncfifo_readable;
wire [9:0] videosoc_uart_tx_fifo_syncfifo_din;
wire [9:0] videosoc_uart_tx_fifo_syncfifo_dout;
reg [4:0] videosoc_uart_tx_fifo_level = 5'd0;
reg videosoc_uart_tx_fifo_replace = 1'd0;
reg [3:0] videosoc_uart_tx_fifo_produce = 4'd0;
reg [3:0] videosoc_uart_tx_fifo_consume = 4'd0;
reg [3:0] videosoc_uart_tx_fifo_wrport_adr = 4'd0;
wire [9:0] videosoc_uart_tx_fifo_wrport_dat_r;
wire videosoc_uart_tx_fifo_wrport_we;
wire [9:0] videosoc_uart_tx_fifo_wrport_dat_w;
wire videosoc_uart_tx_fifo_do_read;
wire [3:0] videosoc_uart_tx_fifo_rdport_adr;
wire [9:0] videosoc_uart_tx_fifo_rdport_dat_r;
wire [7:0] videosoc_uart_tx_fifo_fifo_in_payload_data;
wire videosoc_uart_tx_fifo_fifo_in_first;
wire videosoc_uart_tx_fifo_fifo_in_last;
wire [7:0] videosoc_uart_tx_fifo_fifo_out_payload_data;
wire videosoc_uart_tx_fifo_fifo_out_first;
wire videosoc_uart_tx_fifo_fifo_out_last;
wire videosoc_uart_rx_fifo_sink_valid;
wire videosoc_uart_rx_fifo_sink_ready;
wire videosoc_uart_rx_fifo_sink_first;
wire videosoc_uart_rx_fifo_sink_last;
wire [7:0] videosoc_uart_rx_fifo_sink_payload_data;
wire videosoc_uart_rx_fifo_source_valid;
wire videosoc_uart_rx_fifo_source_ready;
wire videosoc_uart_rx_fifo_source_first;
wire videosoc_uart_rx_fifo_source_last;
wire [7:0] videosoc_uart_rx_fifo_source_payload_data;
wire videosoc_uart_rx_fifo_syncfifo_we;
wire videosoc_uart_rx_fifo_syncfifo_writable;
wire videosoc_uart_rx_fifo_syncfifo_re;
wire videosoc_uart_rx_fifo_syncfifo_readable;
wire [9:0] videosoc_uart_rx_fifo_syncfifo_din;
wire [9:0] videosoc_uart_rx_fifo_syncfifo_dout;
reg [4:0] videosoc_uart_rx_fifo_level = 5'd0;
reg videosoc_uart_rx_fifo_replace = 1'd0;
reg [3:0] videosoc_uart_rx_fifo_produce = 4'd0;
reg [3:0] videosoc_uart_rx_fifo_consume = 4'd0;
reg [3:0] videosoc_uart_rx_fifo_wrport_adr = 4'd0;
wire [9:0] videosoc_uart_rx_fifo_wrport_dat_r;
wire videosoc_uart_rx_fifo_wrport_we;
wire [9:0] videosoc_uart_rx_fifo_wrport_dat_w;
wire videosoc_uart_rx_fifo_do_read;
wire [3:0] videosoc_uart_rx_fifo_rdport_adr;
wire [9:0] videosoc_uart_rx_fifo_rdport_dat_r;
wire [7:0] videosoc_uart_rx_fifo_fifo_in_payload_data;
wire videosoc_uart_rx_fifo_fifo_in_first;
wire videosoc_uart_rx_fifo_fifo_in_last;
wire [7:0] videosoc_uart_rx_fifo_fifo_out_payload_data;
wire videosoc_uart_rx_fifo_fifo_out_first;
wire videosoc_uart_rx_fifo_fifo_out_last;
wire [29:0] videosoc_bridge_wishbone_adr;
wire [31:0] videosoc_bridge_wishbone_dat_w;
wire [31:0] videosoc_bridge_wishbone_dat_r;
wire [3:0] videosoc_bridge_wishbone_sel;
reg videosoc_bridge_wishbone_cyc = 1'd0;
reg videosoc_bridge_wishbone_stb = 1'd0;
wire videosoc_bridge_wishbone_ack;
reg videosoc_bridge_wishbone_we = 1'd0;
reg [2:0] videosoc_bridge_wishbone_cti = 3'd0;
reg [1:0] videosoc_bridge_wishbone_bte = 2'd0;
wire videosoc_bridge_wishbone_err;
reg [2:0] videosoc_bridge_byte_counter = 3'd0;
reg videosoc_bridge_byte_counter_reset = 1'd0;
reg videosoc_bridge_byte_counter_ce = 1'd0;
reg [2:0] videosoc_bridge_word_counter = 3'd0;
reg videosoc_bridge_word_counter_reset = 1'd0;
reg videosoc_bridge_word_counter_ce = 1'd0;
reg [7:0] videosoc_bridge_cmd = 8'd0;
reg videosoc_bridge_cmd_ce = 1'd0;
reg [7:0] videosoc_bridge_length = 8'd0;
reg videosoc_bridge_length_ce = 1'd0;
reg [31:0] videosoc_bridge_address = 32'd0;
reg videosoc_bridge_address_ce = 1'd0;
reg [31:0] videosoc_bridge_data = 32'd0;
reg videosoc_bridge_rx_data_ce = 1'd0;
reg videosoc_bridge_tx_data_ce = 1'd0;
wire videosoc_bridge_reset;
wire videosoc_bridge_wait;
wire videosoc_bridge_done;
reg [23:0] videosoc_bridge_count = 24'd10000000;
reg videosoc_bridge_is_ongoing = 1'd0;
reg [31:0] videosoc_uart_phy_storage_full = 32'd4947802;
wire [31:0] videosoc_uart_phy_storage;
reg videosoc_uart_phy_re = 1'd0;
reg videosoc_uart_phy_sink_valid = 1'd0;
reg videosoc_uart_phy_sink_ready = 1'd0;
reg videosoc_uart_phy_sink_first = 1'd0;
reg videosoc_uart_phy_sink_last = 1'd0;
reg [7:0] videosoc_uart_phy_sink_payload_data = 8'd0;
reg videosoc_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] videosoc_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] videosoc_uart_phy_tx_reg = 8'd0;
reg [3:0] videosoc_uart_phy_tx_bitcount = 4'd0;
reg videosoc_uart_phy_tx_busy = 1'd0;
reg videosoc_uart_phy_source_valid = 1'd0;
reg videosoc_uart_phy_source_ready = 1'd0;
reg videosoc_uart_phy_source_first = 1'd0;
reg videosoc_uart_phy_source_last = 1'd0;
reg [7:0] videosoc_uart_phy_source_payload_data = 8'd0;
reg videosoc_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] videosoc_uart_phy_phase_accumulator_rx = 32'd0;
wire videosoc_uart_phy_rx;
reg videosoc_uart_phy_rx_r = 1'd0;
reg [7:0] videosoc_uart_phy_rx_reg = 8'd0;
reg [3:0] videosoc_uart_phy_rx_bitcount = 4'd0;
reg videosoc_uart_phy_rx_busy = 1'd0;
wire videosoc_sel;
reg [56:0] videosoc_info_dna_status = 57'd0;
wire videosoc_info_dna_do;
reg [6:0] videosoc_info_dna_cnt = 7'd0;
wire [159:0] videosoc_info_git_status;
wire [63:0] videosoc_info_platform_status;
wire [63:0] videosoc_info_target_status;
reg [11:0] videosoc_info_temperature_status = 12'd0;
reg [11:0] videosoc_info_vccint_status = 12'd0;
reg [11:0] videosoc_info_vccaux_status = 12'd0;
reg [11:0] videosoc_info_vccbram_status = 12'd0;
wire [7:0] videosoc_info_alarm;
wire videosoc_info_ot;
wire videosoc_info_busy;
wire [6:0] videosoc_info_channel;
wire videosoc_info_eoc;
wire videosoc_info_eos;
wire [15:0] videosoc_info_data;
wire videosoc_info_drdy;
wire videosoc_oled_spi_pads_cs_n;
reg videosoc_oled_spi_pads_clk = 1'd0;
reg videosoc_oled_spi_pads_mosi = 1'd0;
wire videosoc_oled_spimaster_ctrl_re;
wire videosoc_oled_spimaster_ctrl_r;
reg videosoc_oled_spimaster_ctrl_w = 1'd0;
reg [7:0] videosoc_oled_spimaster_length_storage_full = 8'd0;
wire [7:0] videosoc_oled_spimaster_length_storage;
reg videosoc_oled_spimaster_length_re = 1'd0;
wire videosoc_oled_spimaster_status;
reg [7:0] videosoc_oled_spimaster_mosi_storage_full = 8'd0;
wire [7:0] videosoc_oled_spimaster_mosi_storage;
reg videosoc_oled_spimaster_mosi_re = 1'd0;
reg videosoc_oled_spimaster_irq = 1'd0;
wire videosoc_oled_spimaster_start;
reg videosoc_oled_spimaster_enable_cs = 1'd0;
reg videosoc_oled_spimaster_enable_shift = 1'd0;
reg videosoc_oled_spimaster_done = 1'd0;
reg [3:0] videosoc_oled_spimaster_i = 4'd0;
wire videosoc_oled_spimaster_set_clk;
wire videosoc_oled_spimaster_clr_clk;
reg [7:0] videosoc_oled_spimaster_cnt = 8'd0;
reg videosoc_oled_spimaster_clr_cnt = 1'd0;
reg videosoc_oled_spimaster_inc_cnt = 1'd0;
reg [7:0] videosoc_oled_spimaster_sr_mosi = 8'd0;
reg videosoc_oled_spimaster = 1'd0;
reg [3:0] videosoc_oled_storage_full = 4'd0;
wire [3:0] videosoc_oled_storage;
reg videosoc_oled_re = 1'd0;
reg [1:0] videosoc_ddrphy_storage_full = 2'd0;
wire [1:0] videosoc_ddrphy_storage;
reg videosoc_ddrphy_re = 1'd0;
wire videosoc_ddrphy_rdly_dq_rst_re;
wire videosoc_ddrphy_rdly_dq_rst_r;
reg videosoc_ddrphy_rdly_dq_rst_w = 1'd0;
wire videosoc_ddrphy_rdly_dq_inc_re;
wire videosoc_ddrphy_rdly_dq_inc_r;
reg videosoc_ddrphy_rdly_dq_inc_w = 1'd0;
wire videosoc_ddrphy_rdly_dq_bitslip_re;
wire videosoc_ddrphy_rdly_dq_bitslip_r;
reg videosoc_ddrphy_rdly_dq_bitslip_w = 1'd0;
wire [14:0] videosoc_ddrphy_dfi_p0_address;
wire [2:0] videosoc_ddrphy_dfi_p0_bank;
wire videosoc_ddrphy_dfi_p0_cas_n;
wire videosoc_ddrphy_dfi_p0_cs_n;
wire videosoc_ddrphy_dfi_p0_ras_n;
wire videosoc_ddrphy_dfi_p0_we_n;
wire videosoc_ddrphy_dfi_p0_cke;
wire videosoc_ddrphy_dfi_p0_odt;
wire videosoc_ddrphy_dfi_p0_reset_n;
wire [31:0] videosoc_ddrphy_dfi_p0_wrdata;
wire videosoc_ddrphy_dfi_p0_wrdata_en;
wire [3:0] videosoc_ddrphy_dfi_p0_wrdata_mask;
wire videosoc_ddrphy_dfi_p0_rddata_en;
wire [31:0] videosoc_ddrphy_dfi_p0_rddata;
reg videosoc_ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [14:0] videosoc_ddrphy_dfi_p1_address;
wire [2:0] videosoc_ddrphy_dfi_p1_bank;
wire videosoc_ddrphy_dfi_p1_cas_n;
wire videosoc_ddrphy_dfi_p1_cs_n;
wire videosoc_ddrphy_dfi_p1_ras_n;
wire videosoc_ddrphy_dfi_p1_we_n;
wire videosoc_ddrphy_dfi_p1_cke;
wire videosoc_ddrphy_dfi_p1_odt;
wire videosoc_ddrphy_dfi_p1_reset_n;
wire [31:0] videosoc_ddrphy_dfi_p1_wrdata;
wire videosoc_ddrphy_dfi_p1_wrdata_en;
wire [3:0] videosoc_ddrphy_dfi_p1_wrdata_mask;
wire videosoc_ddrphy_dfi_p1_rddata_en;
wire [31:0] videosoc_ddrphy_dfi_p1_rddata;
reg videosoc_ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [14:0] videosoc_ddrphy_dfi_p2_address;
wire [2:0] videosoc_ddrphy_dfi_p2_bank;
wire videosoc_ddrphy_dfi_p2_cas_n;
wire videosoc_ddrphy_dfi_p2_cs_n;
wire videosoc_ddrphy_dfi_p2_ras_n;
wire videosoc_ddrphy_dfi_p2_we_n;
wire videosoc_ddrphy_dfi_p2_cke;
wire videosoc_ddrphy_dfi_p2_odt;
wire videosoc_ddrphy_dfi_p2_reset_n;
wire [31:0] videosoc_ddrphy_dfi_p2_wrdata;
wire videosoc_ddrphy_dfi_p2_wrdata_en;
wire [3:0] videosoc_ddrphy_dfi_p2_wrdata_mask;
wire videosoc_ddrphy_dfi_p2_rddata_en;
wire [31:0] videosoc_ddrphy_dfi_p2_rddata;
reg videosoc_ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [14:0] videosoc_ddrphy_dfi_p3_address;
wire [2:0] videosoc_ddrphy_dfi_p3_bank;
wire videosoc_ddrphy_dfi_p3_cas_n;
wire videosoc_ddrphy_dfi_p3_cs_n;
wire videosoc_ddrphy_dfi_p3_ras_n;
wire videosoc_ddrphy_dfi_p3_we_n;
wire videosoc_ddrphy_dfi_p3_cke;
wire videosoc_ddrphy_dfi_p3_odt;
wire videosoc_ddrphy_dfi_p3_reset_n;
wire [31:0] videosoc_ddrphy_dfi_p3_wrdata;
wire videosoc_ddrphy_dfi_p3_wrdata_en;
wire [3:0] videosoc_ddrphy_dfi_p3_wrdata_mask;
wire videosoc_ddrphy_dfi_p3_rddata_en;
wire [31:0] videosoc_ddrphy_dfi_p3_rddata;
reg videosoc_ddrphy_dfi_p3_rddata_valid = 1'd0;
wire videosoc_ddrphy_sd_clk_se;
reg videosoc_ddrphy_oe_dqs = 1'd0;
reg [7:0] videosoc_ddrphy_dqs_serdes_pattern = 8'd85;
wire videosoc_ddrphy_dqs0;
wire videosoc_ddrphy_dqs_t0;
wire videosoc_ddrphy_dqs1;
wire videosoc_ddrphy_dqs_t1;
reg videosoc_ddrphy_oe_dq = 1'd0;
wire videosoc_ddrphy_dq_o0;
wire videosoc_ddrphy_dq_i_nodelay0;
wire videosoc_ddrphy_dq_i_delayed0;
wire videosoc_ddrphy_dq_t0;
wire videosoc_ddrphy_dq_o1;
wire videosoc_ddrphy_dq_i_nodelay1;
wire videosoc_ddrphy_dq_i_delayed1;
wire videosoc_ddrphy_dq_t1;
wire videosoc_ddrphy_dq_o2;
wire videosoc_ddrphy_dq_i_nodelay2;
wire videosoc_ddrphy_dq_i_delayed2;
wire videosoc_ddrphy_dq_t2;
wire videosoc_ddrphy_dq_o3;
wire videosoc_ddrphy_dq_i_nodelay3;
wire videosoc_ddrphy_dq_i_delayed3;
wire videosoc_ddrphy_dq_t3;
wire videosoc_ddrphy_dq_o4;
wire videosoc_ddrphy_dq_i_nodelay4;
wire videosoc_ddrphy_dq_i_delayed4;
wire videosoc_ddrphy_dq_t4;
wire videosoc_ddrphy_dq_o5;
wire videosoc_ddrphy_dq_i_nodelay5;
wire videosoc_ddrphy_dq_i_delayed5;
wire videosoc_ddrphy_dq_t5;
wire videosoc_ddrphy_dq_o6;
wire videosoc_ddrphy_dq_i_nodelay6;
wire videosoc_ddrphy_dq_i_delayed6;
wire videosoc_ddrphy_dq_t6;
wire videosoc_ddrphy_dq_o7;
wire videosoc_ddrphy_dq_i_nodelay7;
wire videosoc_ddrphy_dq_i_delayed7;
wire videosoc_ddrphy_dq_t7;
wire videosoc_ddrphy_dq_o8;
wire videosoc_ddrphy_dq_i_nodelay8;
wire videosoc_ddrphy_dq_i_delayed8;
wire videosoc_ddrphy_dq_t8;
wire videosoc_ddrphy_dq_o9;
wire videosoc_ddrphy_dq_i_nodelay9;
wire videosoc_ddrphy_dq_i_delayed9;
wire videosoc_ddrphy_dq_t9;
wire videosoc_ddrphy_dq_o10;
wire videosoc_ddrphy_dq_i_nodelay10;
wire videosoc_ddrphy_dq_i_delayed10;
wire videosoc_ddrphy_dq_t10;
wire videosoc_ddrphy_dq_o11;
wire videosoc_ddrphy_dq_i_nodelay11;
wire videosoc_ddrphy_dq_i_delayed11;
wire videosoc_ddrphy_dq_t11;
wire videosoc_ddrphy_dq_o12;
wire videosoc_ddrphy_dq_i_nodelay12;
wire videosoc_ddrphy_dq_i_delayed12;
wire videosoc_ddrphy_dq_t12;
wire videosoc_ddrphy_dq_o13;
wire videosoc_ddrphy_dq_i_nodelay13;
wire videosoc_ddrphy_dq_i_delayed13;
wire videosoc_ddrphy_dq_t13;
wire videosoc_ddrphy_dq_o14;
wire videosoc_ddrphy_dq_i_nodelay14;
wire videosoc_ddrphy_dq_i_delayed14;
wire videosoc_ddrphy_dq_t14;
wire videosoc_ddrphy_dq_o15;
wire videosoc_ddrphy_dq_i_nodelay15;
wire videosoc_ddrphy_dq_i_delayed15;
wire videosoc_ddrphy_dq_t15;
reg videosoc_ddrphy_n_rddata_en0 = 1'd0;
reg videosoc_ddrphy_n_rddata_en1 = 1'd0;
reg videosoc_ddrphy_n_rddata_en2 = 1'd0;
reg videosoc_ddrphy_n_rddata_en3 = 1'd0;
reg videosoc_ddrphy_n_rddata_en4 = 1'd0;
wire videosoc_ddrphy_oe;
reg [3:0] videosoc_ddrphy_last_wrdata_en = 4'd0;
wire [14:0] videosoc_sdram_inti_p0_address;
wire [2:0] videosoc_sdram_inti_p0_bank;
reg videosoc_sdram_inti_p0_cas_n = 1'd1;
reg videosoc_sdram_inti_p0_cs_n = 1'd1;
reg videosoc_sdram_inti_p0_ras_n = 1'd1;
reg videosoc_sdram_inti_p0_we_n = 1'd1;
wire videosoc_sdram_inti_p0_cke;
wire videosoc_sdram_inti_p0_odt;
wire videosoc_sdram_inti_p0_reset_n;
wire [31:0] videosoc_sdram_inti_p0_wrdata;
wire videosoc_sdram_inti_p0_wrdata_en;
wire [3:0] videosoc_sdram_inti_p0_wrdata_mask;
wire videosoc_sdram_inti_p0_rddata_en;
reg [31:0] videosoc_sdram_inti_p0_rddata = 32'd0;
reg videosoc_sdram_inti_p0_rddata_valid = 1'd0;
wire [14:0] videosoc_sdram_inti_p1_address;
wire [2:0] videosoc_sdram_inti_p1_bank;
reg videosoc_sdram_inti_p1_cas_n = 1'd1;
reg videosoc_sdram_inti_p1_cs_n = 1'd1;
reg videosoc_sdram_inti_p1_ras_n = 1'd1;
reg videosoc_sdram_inti_p1_we_n = 1'd1;
wire videosoc_sdram_inti_p1_cke;
wire videosoc_sdram_inti_p1_odt;
wire videosoc_sdram_inti_p1_reset_n;
wire [31:0] videosoc_sdram_inti_p1_wrdata;
wire videosoc_sdram_inti_p1_wrdata_en;
wire [3:0] videosoc_sdram_inti_p1_wrdata_mask;
wire videosoc_sdram_inti_p1_rddata_en;
reg [31:0] videosoc_sdram_inti_p1_rddata = 32'd0;
reg videosoc_sdram_inti_p1_rddata_valid = 1'd0;
wire [14:0] videosoc_sdram_inti_p2_address;
wire [2:0] videosoc_sdram_inti_p2_bank;
reg videosoc_sdram_inti_p2_cas_n = 1'd1;
reg videosoc_sdram_inti_p2_cs_n = 1'd1;
reg videosoc_sdram_inti_p2_ras_n = 1'd1;
reg videosoc_sdram_inti_p2_we_n = 1'd1;
wire videosoc_sdram_inti_p2_cke;
wire videosoc_sdram_inti_p2_odt;
wire videosoc_sdram_inti_p2_reset_n;
wire [31:0] videosoc_sdram_inti_p2_wrdata;
wire videosoc_sdram_inti_p2_wrdata_en;
wire [3:0] videosoc_sdram_inti_p2_wrdata_mask;
wire videosoc_sdram_inti_p2_rddata_en;
reg [31:0] videosoc_sdram_inti_p2_rddata = 32'd0;
reg videosoc_sdram_inti_p2_rddata_valid = 1'd0;
wire [14:0] videosoc_sdram_inti_p3_address;
wire [2:0] videosoc_sdram_inti_p3_bank;
reg videosoc_sdram_inti_p3_cas_n = 1'd1;
reg videosoc_sdram_inti_p3_cs_n = 1'd1;
reg videosoc_sdram_inti_p3_ras_n = 1'd1;
reg videosoc_sdram_inti_p3_we_n = 1'd1;
wire videosoc_sdram_inti_p3_cke;
wire videosoc_sdram_inti_p3_odt;
wire videosoc_sdram_inti_p3_reset_n;
wire [31:0] videosoc_sdram_inti_p3_wrdata;
wire videosoc_sdram_inti_p3_wrdata_en;
wire [3:0] videosoc_sdram_inti_p3_wrdata_mask;
wire videosoc_sdram_inti_p3_rddata_en;
reg [31:0] videosoc_sdram_inti_p3_rddata = 32'd0;
reg videosoc_sdram_inti_p3_rddata_valid = 1'd0;
wire [14:0] videosoc_sdram_slave_p0_address;
wire [2:0] videosoc_sdram_slave_p0_bank;
wire videosoc_sdram_slave_p0_cas_n;
wire videosoc_sdram_slave_p0_cs_n;
wire videosoc_sdram_slave_p0_ras_n;
wire videosoc_sdram_slave_p0_we_n;
wire videosoc_sdram_slave_p0_cke;
wire videosoc_sdram_slave_p0_odt;
wire videosoc_sdram_slave_p0_reset_n;
wire [31:0] videosoc_sdram_slave_p0_wrdata;
wire videosoc_sdram_slave_p0_wrdata_en;
wire [3:0] videosoc_sdram_slave_p0_wrdata_mask;
wire videosoc_sdram_slave_p0_rddata_en;
reg [31:0] videosoc_sdram_slave_p0_rddata = 32'd0;
reg videosoc_sdram_slave_p0_rddata_valid = 1'd0;
wire [14:0] videosoc_sdram_slave_p1_address;
wire [2:0] videosoc_sdram_slave_p1_bank;
wire videosoc_sdram_slave_p1_cas_n;
wire videosoc_sdram_slave_p1_cs_n;
wire videosoc_sdram_slave_p1_ras_n;
wire videosoc_sdram_slave_p1_we_n;
wire videosoc_sdram_slave_p1_cke;
wire videosoc_sdram_slave_p1_odt;
wire videosoc_sdram_slave_p1_reset_n;
wire [31:0] videosoc_sdram_slave_p1_wrdata;
wire videosoc_sdram_slave_p1_wrdata_en;
wire [3:0] videosoc_sdram_slave_p1_wrdata_mask;
wire videosoc_sdram_slave_p1_rddata_en;
reg [31:0] videosoc_sdram_slave_p1_rddata = 32'd0;
reg videosoc_sdram_slave_p1_rddata_valid = 1'd0;
wire [14:0] videosoc_sdram_slave_p2_address;
wire [2:0] videosoc_sdram_slave_p2_bank;
wire videosoc_sdram_slave_p2_cas_n;
wire videosoc_sdram_slave_p2_cs_n;
wire videosoc_sdram_slave_p2_ras_n;
wire videosoc_sdram_slave_p2_we_n;
wire videosoc_sdram_slave_p2_cke;
wire videosoc_sdram_slave_p2_odt;
wire videosoc_sdram_slave_p2_reset_n;
wire [31:0] videosoc_sdram_slave_p2_wrdata;
wire videosoc_sdram_slave_p2_wrdata_en;
wire [3:0] videosoc_sdram_slave_p2_wrdata_mask;
wire videosoc_sdram_slave_p2_rddata_en;
reg [31:0] videosoc_sdram_slave_p2_rddata = 32'd0;
reg videosoc_sdram_slave_p2_rddata_valid = 1'd0;
wire [14:0] videosoc_sdram_slave_p3_address;
wire [2:0] videosoc_sdram_slave_p3_bank;
wire videosoc_sdram_slave_p3_cas_n;
wire videosoc_sdram_slave_p3_cs_n;
wire videosoc_sdram_slave_p3_ras_n;
wire videosoc_sdram_slave_p3_we_n;
wire videosoc_sdram_slave_p3_cke;
wire videosoc_sdram_slave_p3_odt;
wire videosoc_sdram_slave_p3_reset_n;
wire [31:0] videosoc_sdram_slave_p3_wrdata;
wire videosoc_sdram_slave_p3_wrdata_en;
wire [3:0] videosoc_sdram_slave_p3_wrdata_mask;
wire videosoc_sdram_slave_p3_rddata_en;
reg [31:0] videosoc_sdram_slave_p3_rddata = 32'd0;
reg videosoc_sdram_slave_p3_rddata_valid = 1'd0;
reg [14:0] videosoc_sdram_master_p0_address = 15'd0;
reg [2:0] videosoc_sdram_master_p0_bank = 3'd0;
reg videosoc_sdram_master_p0_cas_n = 1'd1;
reg videosoc_sdram_master_p0_cs_n = 1'd1;
reg videosoc_sdram_master_p0_ras_n = 1'd1;
reg videosoc_sdram_master_p0_we_n = 1'd1;
reg videosoc_sdram_master_p0_cke = 1'd0;
reg videosoc_sdram_master_p0_odt = 1'd0;
reg videosoc_sdram_master_p0_reset_n = 1'd0;
reg [31:0] videosoc_sdram_master_p0_wrdata = 32'd0;
reg videosoc_sdram_master_p0_wrdata_en = 1'd0;
reg [3:0] videosoc_sdram_master_p0_wrdata_mask = 4'd0;
reg videosoc_sdram_master_p0_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_master_p0_rddata;
wire videosoc_sdram_master_p0_rddata_valid;
reg [14:0] videosoc_sdram_master_p1_address = 15'd0;
reg [2:0] videosoc_sdram_master_p1_bank = 3'd0;
reg videosoc_sdram_master_p1_cas_n = 1'd1;
reg videosoc_sdram_master_p1_cs_n = 1'd1;
reg videosoc_sdram_master_p1_ras_n = 1'd1;
reg videosoc_sdram_master_p1_we_n = 1'd1;
reg videosoc_sdram_master_p1_cke = 1'd0;
reg videosoc_sdram_master_p1_odt = 1'd0;
reg videosoc_sdram_master_p1_reset_n = 1'd0;
reg [31:0] videosoc_sdram_master_p1_wrdata = 32'd0;
reg videosoc_sdram_master_p1_wrdata_en = 1'd0;
reg [3:0] videosoc_sdram_master_p1_wrdata_mask = 4'd0;
reg videosoc_sdram_master_p1_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_master_p1_rddata;
wire videosoc_sdram_master_p1_rddata_valid;
reg [14:0] videosoc_sdram_master_p2_address = 15'd0;
reg [2:0] videosoc_sdram_master_p2_bank = 3'd0;
reg videosoc_sdram_master_p2_cas_n = 1'd1;
reg videosoc_sdram_master_p2_cs_n = 1'd1;
reg videosoc_sdram_master_p2_ras_n = 1'd1;
reg videosoc_sdram_master_p2_we_n = 1'd1;
reg videosoc_sdram_master_p2_cke = 1'd0;
reg videosoc_sdram_master_p2_odt = 1'd0;
reg videosoc_sdram_master_p2_reset_n = 1'd0;
reg [31:0] videosoc_sdram_master_p2_wrdata = 32'd0;
reg videosoc_sdram_master_p2_wrdata_en = 1'd0;
reg [3:0] videosoc_sdram_master_p2_wrdata_mask = 4'd0;
reg videosoc_sdram_master_p2_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_master_p2_rddata;
wire videosoc_sdram_master_p2_rddata_valid;
reg [14:0] videosoc_sdram_master_p3_address = 15'd0;
reg [2:0] videosoc_sdram_master_p3_bank = 3'd0;
reg videosoc_sdram_master_p3_cas_n = 1'd1;
reg videosoc_sdram_master_p3_cs_n = 1'd1;
reg videosoc_sdram_master_p3_ras_n = 1'd1;
reg videosoc_sdram_master_p3_we_n = 1'd1;
reg videosoc_sdram_master_p3_cke = 1'd0;
reg videosoc_sdram_master_p3_odt = 1'd0;
reg videosoc_sdram_master_p3_reset_n = 1'd0;
reg [31:0] videosoc_sdram_master_p3_wrdata = 32'd0;
reg videosoc_sdram_master_p3_wrdata_en = 1'd0;
reg [3:0] videosoc_sdram_master_p3_wrdata_mask = 4'd0;
reg videosoc_sdram_master_p3_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_master_p3_rddata;
wire videosoc_sdram_master_p3_rddata_valid;
reg [3:0] videosoc_sdram_storage_full = 4'd0;
wire [3:0] videosoc_sdram_storage;
reg videosoc_sdram_re = 1'd0;
reg [5:0] videosoc_sdram_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] videosoc_sdram_phaseinjector0_command_storage;
reg videosoc_sdram_phaseinjector0_command_re = 1'd0;
wire videosoc_sdram_phaseinjector0_command_issue_re;
wire videosoc_sdram_phaseinjector0_command_issue_r;
reg videosoc_sdram_phaseinjector0_command_issue_w = 1'd0;
reg [14:0] videosoc_sdram_phaseinjector0_address_storage_full = 15'd0;
wire [14:0] videosoc_sdram_phaseinjector0_address_storage;
reg videosoc_sdram_phaseinjector0_address_re = 1'd0;
reg [2:0] videosoc_sdram_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] videosoc_sdram_phaseinjector0_baddress_storage;
reg videosoc_sdram_phaseinjector0_baddress_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector0_wrdata_storage_full = 32'd0;
wire [31:0] videosoc_sdram_phaseinjector0_wrdata_storage;
reg videosoc_sdram_phaseinjector0_wrdata_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector0_status = 32'd0;
reg [5:0] videosoc_sdram_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] videosoc_sdram_phaseinjector1_command_storage;
reg videosoc_sdram_phaseinjector1_command_re = 1'd0;
wire videosoc_sdram_phaseinjector1_command_issue_re;
wire videosoc_sdram_phaseinjector1_command_issue_r;
reg videosoc_sdram_phaseinjector1_command_issue_w = 1'd0;
reg [14:0] videosoc_sdram_phaseinjector1_address_storage_full = 15'd0;
wire [14:0] videosoc_sdram_phaseinjector1_address_storage;
reg videosoc_sdram_phaseinjector1_address_re = 1'd0;
reg [2:0] videosoc_sdram_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] videosoc_sdram_phaseinjector1_baddress_storage;
reg videosoc_sdram_phaseinjector1_baddress_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector1_wrdata_storage_full = 32'd0;
wire [31:0] videosoc_sdram_phaseinjector1_wrdata_storage;
reg videosoc_sdram_phaseinjector1_wrdata_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector1_status = 32'd0;
reg [5:0] videosoc_sdram_phaseinjector2_command_storage_full = 6'd0;
wire [5:0] videosoc_sdram_phaseinjector2_command_storage;
reg videosoc_sdram_phaseinjector2_command_re = 1'd0;
wire videosoc_sdram_phaseinjector2_command_issue_re;
wire videosoc_sdram_phaseinjector2_command_issue_r;
reg videosoc_sdram_phaseinjector2_command_issue_w = 1'd0;
reg [14:0] videosoc_sdram_phaseinjector2_address_storage_full = 15'd0;
wire [14:0] videosoc_sdram_phaseinjector2_address_storage;
reg videosoc_sdram_phaseinjector2_address_re = 1'd0;
reg [2:0] videosoc_sdram_phaseinjector2_baddress_storage_full = 3'd0;
wire [2:0] videosoc_sdram_phaseinjector2_baddress_storage;
reg videosoc_sdram_phaseinjector2_baddress_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector2_wrdata_storage_full = 32'd0;
wire [31:0] videosoc_sdram_phaseinjector2_wrdata_storage;
reg videosoc_sdram_phaseinjector2_wrdata_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector2_status = 32'd0;
reg [5:0] videosoc_sdram_phaseinjector3_command_storage_full = 6'd0;
wire [5:0] videosoc_sdram_phaseinjector3_command_storage;
reg videosoc_sdram_phaseinjector3_command_re = 1'd0;
wire videosoc_sdram_phaseinjector3_command_issue_re;
wire videosoc_sdram_phaseinjector3_command_issue_r;
reg videosoc_sdram_phaseinjector3_command_issue_w = 1'd0;
reg [14:0] videosoc_sdram_phaseinjector3_address_storage_full = 15'd0;
wire [14:0] videosoc_sdram_phaseinjector3_address_storage;
reg videosoc_sdram_phaseinjector3_address_re = 1'd0;
reg [2:0] videosoc_sdram_phaseinjector3_baddress_storage_full = 3'd0;
wire [2:0] videosoc_sdram_phaseinjector3_baddress_storage;
reg videosoc_sdram_phaseinjector3_baddress_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector3_wrdata_storage_full = 32'd0;
wire [31:0] videosoc_sdram_phaseinjector3_wrdata_storage;
reg videosoc_sdram_phaseinjector3_wrdata_re = 1'd0;
reg [31:0] videosoc_sdram_phaseinjector3_status = 32'd0;
reg [14:0] videosoc_sdram_dfi_p0_address = 15'd0;
reg [2:0] videosoc_sdram_dfi_p0_bank = 3'd0;
reg videosoc_sdram_dfi_p0_cas_n = 1'd1;
wire videosoc_sdram_dfi_p0_cs_n;
reg videosoc_sdram_dfi_p0_ras_n = 1'd1;
reg videosoc_sdram_dfi_p0_we_n = 1'd1;
wire videosoc_sdram_dfi_p0_cke;
wire videosoc_sdram_dfi_p0_odt;
wire videosoc_sdram_dfi_p0_reset_n;
wire [31:0] videosoc_sdram_dfi_p0_wrdata;
reg videosoc_sdram_dfi_p0_wrdata_en = 1'd0;
wire [3:0] videosoc_sdram_dfi_p0_wrdata_mask;
reg videosoc_sdram_dfi_p0_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_dfi_p0_rddata;
wire videosoc_sdram_dfi_p0_rddata_valid;
reg [14:0] videosoc_sdram_dfi_p1_address = 15'd0;
reg [2:0] videosoc_sdram_dfi_p1_bank = 3'd0;
reg videosoc_sdram_dfi_p1_cas_n = 1'd1;
wire videosoc_sdram_dfi_p1_cs_n;
reg videosoc_sdram_dfi_p1_ras_n = 1'd1;
reg videosoc_sdram_dfi_p1_we_n = 1'd1;
wire videosoc_sdram_dfi_p1_cke;
wire videosoc_sdram_dfi_p1_odt;
wire videosoc_sdram_dfi_p1_reset_n;
wire [31:0] videosoc_sdram_dfi_p1_wrdata;
reg videosoc_sdram_dfi_p1_wrdata_en = 1'd0;
wire [3:0] videosoc_sdram_dfi_p1_wrdata_mask;
reg videosoc_sdram_dfi_p1_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_dfi_p1_rddata;
wire videosoc_sdram_dfi_p1_rddata_valid;
reg [14:0] videosoc_sdram_dfi_p2_address = 15'd0;
reg [2:0] videosoc_sdram_dfi_p2_bank = 3'd0;
reg videosoc_sdram_dfi_p2_cas_n = 1'd1;
wire videosoc_sdram_dfi_p2_cs_n;
reg videosoc_sdram_dfi_p2_ras_n = 1'd1;
reg videosoc_sdram_dfi_p2_we_n = 1'd1;
wire videosoc_sdram_dfi_p2_cke;
wire videosoc_sdram_dfi_p2_odt;
wire videosoc_sdram_dfi_p2_reset_n;
wire [31:0] videosoc_sdram_dfi_p2_wrdata;
reg videosoc_sdram_dfi_p2_wrdata_en = 1'd0;
wire [3:0] videosoc_sdram_dfi_p2_wrdata_mask;
reg videosoc_sdram_dfi_p2_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_dfi_p2_rddata;
wire videosoc_sdram_dfi_p2_rddata_valid;
reg [14:0] videosoc_sdram_dfi_p3_address = 15'd0;
reg [2:0] videosoc_sdram_dfi_p3_bank = 3'd0;
reg videosoc_sdram_dfi_p3_cas_n = 1'd1;
wire videosoc_sdram_dfi_p3_cs_n;
reg videosoc_sdram_dfi_p3_ras_n = 1'd1;
reg videosoc_sdram_dfi_p3_we_n = 1'd1;
wire videosoc_sdram_dfi_p3_cke;
wire videosoc_sdram_dfi_p3_odt;
wire videosoc_sdram_dfi_p3_reset_n;
wire [31:0] videosoc_sdram_dfi_p3_wrdata;
reg videosoc_sdram_dfi_p3_wrdata_en = 1'd0;
wire [3:0] videosoc_sdram_dfi_p3_wrdata_mask;
reg videosoc_sdram_dfi_p3_rddata_en = 1'd0;
wire [31:0] videosoc_sdram_dfi_p3_rddata;
wire videosoc_sdram_dfi_p3_rddata_valid;
wire videosoc_sdram_interface_bank0_valid;
wire videosoc_sdram_interface_bank0_ready;
wire videosoc_sdram_interface_bank0_we;
wire [21:0] videosoc_sdram_interface_bank0_adr;
wire videosoc_sdram_interface_bank0_lock;
wire videosoc_sdram_interface_bank0_wdata_ready;
wire videosoc_sdram_interface_bank0_rdata_valid;
wire videosoc_sdram_interface_bank1_valid;
wire videosoc_sdram_interface_bank1_ready;
wire videosoc_sdram_interface_bank1_we;
wire [21:0] videosoc_sdram_interface_bank1_adr;
wire videosoc_sdram_interface_bank1_lock;
wire videosoc_sdram_interface_bank1_wdata_ready;
wire videosoc_sdram_interface_bank1_rdata_valid;
wire videosoc_sdram_interface_bank2_valid;
wire videosoc_sdram_interface_bank2_ready;
wire videosoc_sdram_interface_bank2_we;
wire [21:0] videosoc_sdram_interface_bank2_adr;
wire videosoc_sdram_interface_bank2_lock;
wire videosoc_sdram_interface_bank2_wdata_ready;
wire videosoc_sdram_interface_bank2_rdata_valid;
wire videosoc_sdram_interface_bank3_valid;
wire videosoc_sdram_interface_bank3_ready;
wire videosoc_sdram_interface_bank3_we;
wire [21:0] videosoc_sdram_interface_bank3_adr;
wire videosoc_sdram_interface_bank3_lock;
wire videosoc_sdram_interface_bank3_wdata_ready;
wire videosoc_sdram_interface_bank3_rdata_valid;
wire videosoc_sdram_interface_bank4_valid;
wire videosoc_sdram_interface_bank4_ready;
wire videosoc_sdram_interface_bank4_we;
wire [21:0] videosoc_sdram_interface_bank4_adr;
wire videosoc_sdram_interface_bank4_lock;
wire videosoc_sdram_interface_bank4_wdata_ready;
wire videosoc_sdram_interface_bank4_rdata_valid;
wire videosoc_sdram_interface_bank5_valid;
wire videosoc_sdram_interface_bank5_ready;
wire videosoc_sdram_interface_bank5_we;
wire [21:0] videosoc_sdram_interface_bank5_adr;
wire videosoc_sdram_interface_bank5_lock;
wire videosoc_sdram_interface_bank5_wdata_ready;
wire videosoc_sdram_interface_bank5_rdata_valid;
wire videosoc_sdram_interface_bank6_valid;
wire videosoc_sdram_interface_bank6_ready;
wire videosoc_sdram_interface_bank6_we;
wire [21:0] videosoc_sdram_interface_bank6_adr;
wire videosoc_sdram_interface_bank6_lock;
wire videosoc_sdram_interface_bank6_wdata_ready;
wire videosoc_sdram_interface_bank6_rdata_valid;
wire videosoc_sdram_interface_bank7_valid;
wire videosoc_sdram_interface_bank7_ready;
wire videosoc_sdram_interface_bank7_we;
wire [21:0] videosoc_sdram_interface_bank7_adr;
wire videosoc_sdram_interface_bank7_lock;
wire videosoc_sdram_interface_bank7_wdata_ready;
wire videosoc_sdram_interface_bank7_rdata_valid;
reg [127:0] videosoc_sdram_interface_wdata = 128'd0;
reg [15:0] videosoc_sdram_interface_wdata_we = 16'd0;
wire [127:0] videosoc_sdram_interface_rdata;
reg videosoc_sdram_cmd_valid = 1'd0;
reg videosoc_sdram_cmd_ready = 1'd0;
reg videosoc_sdram_cmd_last = 1'd0;
reg [14:0] videosoc_sdram_cmd_payload_a = 15'd0;
reg [2:0] videosoc_sdram_cmd_payload_ba = 3'd0;
reg videosoc_sdram_cmd_payload_cas = 1'd0;
reg videosoc_sdram_cmd_payload_ras = 1'd0;
reg videosoc_sdram_cmd_payload_we = 1'd0;
reg videosoc_sdram_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_cmd_payload_is_write = 1'd0;
reg videosoc_sdram_seq_start = 1'd0;
reg videosoc_sdram_seq_done = 1'd0;
reg [4:0] videosoc_sdram_counter = 5'd0;
wire videosoc_sdram_wait;
wire videosoc_sdram_done;
reg [9:0] videosoc_sdram_count = 10'd782;
wire videosoc_sdram_bankmachine0_req_valid;
wire videosoc_sdram_bankmachine0_req_ready;
wire videosoc_sdram_bankmachine0_req_we;
wire [21:0] videosoc_sdram_bankmachine0_req_adr;
wire videosoc_sdram_bankmachine0_req_lock;
reg videosoc_sdram_bankmachine0_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine0_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine0_refresh_req;
reg videosoc_sdram_bankmachine0_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine0_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine0_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine0_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine0_cmd_payload_ba;
reg videosoc_sdram_bankmachine0_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine0_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine0_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine0_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine0_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine0_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine0_sink_valid;
wire videosoc_sdram_bankmachine0_sink_ready;
reg videosoc_sdram_bankmachine0_sink_first = 1'd0;
reg videosoc_sdram_bankmachine0_sink_last = 1'd0;
wire videosoc_sdram_bankmachine0_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine0_sink_payload_adr;
wire videosoc_sdram_bankmachine0_source_valid;
wire videosoc_sdram_bankmachine0_source_ready;
wire videosoc_sdram_bankmachine0_source_first;
wire videosoc_sdram_bankmachine0_source_last;
wire videosoc_sdram_bankmachine0_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine0_source_payload_adr;
wire videosoc_sdram_bankmachine0_syncfifo0_we;
wire videosoc_sdram_bankmachine0_syncfifo0_writable;
wire videosoc_sdram_bankmachine0_syncfifo0_re;
wire videosoc_sdram_bankmachine0_syncfifo0_readable;
wire [24:0] videosoc_sdram_bankmachine0_syncfifo0_din;
wire [24:0] videosoc_sdram_bankmachine0_syncfifo0_dout;
reg [3:0] videosoc_sdram_bankmachine0_level = 4'd0;
reg videosoc_sdram_bankmachine0_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine0_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine0_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine0_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine0_wrport_dat_r;
wire videosoc_sdram_bankmachine0_wrport_we;
wire [24:0] videosoc_sdram_bankmachine0_wrport_dat_w;
wire videosoc_sdram_bankmachine0_do_read;
wire [2:0] videosoc_sdram_bankmachine0_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine0_rdport_dat_r;
wire videosoc_sdram_bankmachine0_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine0_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine0_fifo_in_first;
wire videosoc_sdram_bankmachine0_fifo_in_last;
wire videosoc_sdram_bankmachine0_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine0_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine0_fifo_out_first;
wire videosoc_sdram_bankmachine0_fifo_out_last;
reg videosoc_sdram_bankmachine0_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine0_openrow = 15'd0;
wire videosoc_sdram_bankmachine0_hit;
reg videosoc_sdram_bankmachine0_track_open = 1'd0;
reg videosoc_sdram_bankmachine0_track_close = 1'd0;
reg videosoc_sdram_bankmachine0_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine0_wait;
wire videosoc_sdram_bankmachine0_done;
reg [2:0] videosoc_sdram_bankmachine0_count = 3'd5;
wire videosoc_sdram_bankmachine1_req_valid;
wire videosoc_sdram_bankmachine1_req_ready;
wire videosoc_sdram_bankmachine1_req_we;
wire [21:0] videosoc_sdram_bankmachine1_req_adr;
wire videosoc_sdram_bankmachine1_req_lock;
reg videosoc_sdram_bankmachine1_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine1_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine1_refresh_req;
reg videosoc_sdram_bankmachine1_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine1_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine1_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine1_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine1_cmd_payload_ba;
reg videosoc_sdram_bankmachine1_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine1_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine1_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine1_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine1_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine1_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine1_sink_valid;
wire videosoc_sdram_bankmachine1_sink_ready;
reg videosoc_sdram_bankmachine1_sink_first = 1'd0;
reg videosoc_sdram_bankmachine1_sink_last = 1'd0;
wire videosoc_sdram_bankmachine1_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine1_sink_payload_adr;
wire videosoc_sdram_bankmachine1_source_valid;
wire videosoc_sdram_bankmachine1_source_ready;
wire videosoc_sdram_bankmachine1_source_first;
wire videosoc_sdram_bankmachine1_source_last;
wire videosoc_sdram_bankmachine1_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine1_source_payload_adr;
wire videosoc_sdram_bankmachine1_syncfifo1_we;
wire videosoc_sdram_bankmachine1_syncfifo1_writable;
wire videosoc_sdram_bankmachine1_syncfifo1_re;
wire videosoc_sdram_bankmachine1_syncfifo1_readable;
wire [24:0] videosoc_sdram_bankmachine1_syncfifo1_din;
wire [24:0] videosoc_sdram_bankmachine1_syncfifo1_dout;
reg [3:0] videosoc_sdram_bankmachine1_level = 4'd0;
reg videosoc_sdram_bankmachine1_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine1_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine1_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine1_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine1_wrport_dat_r;
wire videosoc_sdram_bankmachine1_wrport_we;
wire [24:0] videosoc_sdram_bankmachine1_wrport_dat_w;
wire videosoc_sdram_bankmachine1_do_read;
wire [2:0] videosoc_sdram_bankmachine1_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine1_rdport_dat_r;
wire videosoc_sdram_bankmachine1_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine1_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine1_fifo_in_first;
wire videosoc_sdram_bankmachine1_fifo_in_last;
wire videosoc_sdram_bankmachine1_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine1_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine1_fifo_out_first;
wire videosoc_sdram_bankmachine1_fifo_out_last;
reg videosoc_sdram_bankmachine1_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine1_openrow = 15'd0;
wire videosoc_sdram_bankmachine1_hit;
reg videosoc_sdram_bankmachine1_track_open = 1'd0;
reg videosoc_sdram_bankmachine1_track_close = 1'd0;
reg videosoc_sdram_bankmachine1_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine1_wait;
wire videosoc_sdram_bankmachine1_done;
reg [2:0] videosoc_sdram_bankmachine1_count = 3'd5;
wire videosoc_sdram_bankmachine2_req_valid;
wire videosoc_sdram_bankmachine2_req_ready;
wire videosoc_sdram_bankmachine2_req_we;
wire [21:0] videosoc_sdram_bankmachine2_req_adr;
wire videosoc_sdram_bankmachine2_req_lock;
reg videosoc_sdram_bankmachine2_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine2_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine2_refresh_req;
reg videosoc_sdram_bankmachine2_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine2_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine2_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine2_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine2_cmd_payload_ba;
reg videosoc_sdram_bankmachine2_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine2_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine2_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine2_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine2_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine2_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine2_sink_valid;
wire videosoc_sdram_bankmachine2_sink_ready;
reg videosoc_sdram_bankmachine2_sink_first = 1'd0;
reg videosoc_sdram_bankmachine2_sink_last = 1'd0;
wire videosoc_sdram_bankmachine2_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine2_sink_payload_adr;
wire videosoc_sdram_bankmachine2_source_valid;
wire videosoc_sdram_bankmachine2_source_ready;
wire videosoc_sdram_bankmachine2_source_first;
wire videosoc_sdram_bankmachine2_source_last;
wire videosoc_sdram_bankmachine2_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine2_source_payload_adr;
wire videosoc_sdram_bankmachine2_syncfifo2_we;
wire videosoc_sdram_bankmachine2_syncfifo2_writable;
wire videosoc_sdram_bankmachine2_syncfifo2_re;
wire videosoc_sdram_bankmachine2_syncfifo2_readable;
wire [24:0] videosoc_sdram_bankmachine2_syncfifo2_din;
wire [24:0] videosoc_sdram_bankmachine2_syncfifo2_dout;
reg [3:0] videosoc_sdram_bankmachine2_level = 4'd0;
reg videosoc_sdram_bankmachine2_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine2_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine2_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine2_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine2_wrport_dat_r;
wire videosoc_sdram_bankmachine2_wrport_we;
wire [24:0] videosoc_sdram_bankmachine2_wrport_dat_w;
wire videosoc_sdram_bankmachine2_do_read;
wire [2:0] videosoc_sdram_bankmachine2_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine2_rdport_dat_r;
wire videosoc_sdram_bankmachine2_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine2_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine2_fifo_in_first;
wire videosoc_sdram_bankmachine2_fifo_in_last;
wire videosoc_sdram_bankmachine2_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine2_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine2_fifo_out_first;
wire videosoc_sdram_bankmachine2_fifo_out_last;
reg videosoc_sdram_bankmachine2_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine2_openrow = 15'd0;
wire videosoc_sdram_bankmachine2_hit;
reg videosoc_sdram_bankmachine2_track_open = 1'd0;
reg videosoc_sdram_bankmachine2_track_close = 1'd0;
reg videosoc_sdram_bankmachine2_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine2_wait;
wire videosoc_sdram_bankmachine2_done;
reg [2:0] videosoc_sdram_bankmachine2_count = 3'd5;
wire videosoc_sdram_bankmachine3_req_valid;
wire videosoc_sdram_bankmachine3_req_ready;
wire videosoc_sdram_bankmachine3_req_we;
wire [21:0] videosoc_sdram_bankmachine3_req_adr;
wire videosoc_sdram_bankmachine3_req_lock;
reg videosoc_sdram_bankmachine3_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine3_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine3_refresh_req;
reg videosoc_sdram_bankmachine3_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine3_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine3_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine3_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine3_cmd_payload_ba;
reg videosoc_sdram_bankmachine3_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine3_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine3_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine3_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine3_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine3_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine3_sink_valid;
wire videosoc_sdram_bankmachine3_sink_ready;
reg videosoc_sdram_bankmachine3_sink_first = 1'd0;
reg videosoc_sdram_bankmachine3_sink_last = 1'd0;
wire videosoc_sdram_bankmachine3_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine3_sink_payload_adr;
wire videosoc_sdram_bankmachine3_source_valid;
wire videosoc_sdram_bankmachine3_source_ready;
wire videosoc_sdram_bankmachine3_source_first;
wire videosoc_sdram_bankmachine3_source_last;
wire videosoc_sdram_bankmachine3_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine3_source_payload_adr;
wire videosoc_sdram_bankmachine3_syncfifo3_we;
wire videosoc_sdram_bankmachine3_syncfifo3_writable;
wire videosoc_sdram_bankmachine3_syncfifo3_re;
wire videosoc_sdram_bankmachine3_syncfifo3_readable;
wire [24:0] videosoc_sdram_bankmachine3_syncfifo3_din;
wire [24:0] videosoc_sdram_bankmachine3_syncfifo3_dout;
reg [3:0] videosoc_sdram_bankmachine3_level = 4'd0;
reg videosoc_sdram_bankmachine3_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine3_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine3_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine3_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine3_wrport_dat_r;
wire videosoc_sdram_bankmachine3_wrport_we;
wire [24:0] videosoc_sdram_bankmachine3_wrport_dat_w;
wire videosoc_sdram_bankmachine3_do_read;
wire [2:0] videosoc_sdram_bankmachine3_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine3_rdport_dat_r;
wire videosoc_sdram_bankmachine3_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine3_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine3_fifo_in_first;
wire videosoc_sdram_bankmachine3_fifo_in_last;
wire videosoc_sdram_bankmachine3_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine3_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine3_fifo_out_first;
wire videosoc_sdram_bankmachine3_fifo_out_last;
reg videosoc_sdram_bankmachine3_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine3_openrow = 15'd0;
wire videosoc_sdram_bankmachine3_hit;
reg videosoc_sdram_bankmachine3_track_open = 1'd0;
reg videosoc_sdram_bankmachine3_track_close = 1'd0;
reg videosoc_sdram_bankmachine3_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine3_wait;
wire videosoc_sdram_bankmachine3_done;
reg [2:0] videosoc_sdram_bankmachine3_count = 3'd5;
wire videosoc_sdram_bankmachine4_req_valid;
wire videosoc_sdram_bankmachine4_req_ready;
wire videosoc_sdram_bankmachine4_req_we;
wire [21:0] videosoc_sdram_bankmachine4_req_adr;
wire videosoc_sdram_bankmachine4_req_lock;
reg videosoc_sdram_bankmachine4_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine4_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine4_refresh_req;
reg videosoc_sdram_bankmachine4_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine4_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine4_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine4_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine4_cmd_payload_ba;
reg videosoc_sdram_bankmachine4_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine4_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine4_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine4_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine4_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine4_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine4_sink_valid;
wire videosoc_sdram_bankmachine4_sink_ready;
reg videosoc_sdram_bankmachine4_sink_first = 1'd0;
reg videosoc_sdram_bankmachine4_sink_last = 1'd0;
wire videosoc_sdram_bankmachine4_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine4_sink_payload_adr;
wire videosoc_sdram_bankmachine4_source_valid;
wire videosoc_sdram_bankmachine4_source_ready;
wire videosoc_sdram_bankmachine4_source_first;
wire videosoc_sdram_bankmachine4_source_last;
wire videosoc_sdram_bankmachine4_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine4_source_payload_adr;
wire videosoc_sdram_bankmachine4_syncfifo4_we;
wire videosoc_sdram_bankmachine4_syncfifo4_writable;
wire videosoc_sdram_bankmachine4_syncfifo4_re;
wire videosoc_sdram_bankmachine4_syncfifo4_readable;
wire [24:0] videosoc_sdram_bankmachine4_syncfifo4_din;
wire [24:0] videosoc_sdram_bankmachine4_syncfifo4_dout;
reg [3:0] videosoc_sdram_bankmachine4_level = 4'd0;
reg videosoc_sdram_bankmachine4_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine4_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine4_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine4_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine4_wrport_dat_r;
wire videosoc_sdram_bankmachine4_wrport_we;
wire [24:0] videosoc_sdram_bankmachine4_wrport_dat_w;
wire videosoc_sdram_bankmachine4_do_read;
wire [2:0] videosoc_sdram_bankmachine4_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine4_rdport_dat_r;
wire videosoc_sdram_bankmachine4_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine4_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine4_fifo_in_first;
wire videosoc_sdram_bankmachine4_fifo_in_last;
wire videosoc_sdram_bankmachine4_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine4_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine4_fifo_out_first;
wire videosoc_sdram_bankmachine4_fifo_out_last;
reg videosoc_sdram_bankmachine4_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine4_openrow = 15'd0;
wire videosoc_sdram_bankmachine4_hit;
reg videosoc_sdram_bankmachine4_track_open = 1'd0;
reg videosoc_sdram_bankmachine4_track_close = 1'd0;
reg videosoc_sdram_bankmachine4_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine4_wait;
wire videosoc_sdram_bankmachine4_done;
reg [2:0] videosoc_sdram_bankmachine4_count = 3'd5;
wire videosoc_sdram_bankmachine5_req_valid;
wire videosoc_sdram_bankmachine5_req_ready;
wire videosoc_sdram_bankmachine5_req_we;
wire [21:0] videosoc_sdram_bankmachine5_req_adr;
wire videosoc_sdram_bankmachine5_req_lock;
reg videosoc_sdram_bankmachine5_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine5_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine5_refresh_req;
reg videosoc_sdram_bankmachine5_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine5_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine5_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine5_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine5_cmd_payload_ba;
reg videosoc_sdram_bankmachine5_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine5_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine5_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine5_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine5_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine5_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine5_sink_valid;
wire videosoc_sdram_bankmachine5_sink_ready;
reg videosoc_sdram_bankmachine5_sink_first = 1'd0;
reg videosoc_sdram_bankmachine5_sink_last = 1'd0;
wire videosoc_sdram_bankmachine5_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine5_sink_payload_adr;
wire videosoc_sdram_bankmachine5_source_valid;
wire videosoc_sdram_bankmachine5_source_ready;
wire videosoc_sdram_bankmachine5_source_first;
wire videosoc_sdram_bankmachine5_source_last;
wire videosoc_sdram_bankmachine5_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine5_source_payload_adr;
wire videosoc_sdram_bankmachine5_syncfifo5_we;
wire videosoc_sdram_bankmachine5_syncfifo5_writable;
wire videosoc_sdram_bankmachine5_syncfifo5_re;
wire videosoc_sdram_bankmachine5_syncfifo5_readable;
wire [24:0] videosoc_sdram_bankmachine5_syncfifo5_din;
wire [24:0] videosoc_sdram_bankmachine5_syncfifo5_dout;
reg [3:0] videosoc_sdram_bankmachine5_level = 4'd0;
reg videosoc_sdram_bankmachine5_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine5_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine5_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine5_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine5_wrport_dat_r;
wire videosoc_sdram_bankmachine5_wrport_we;
wire [24:0] videosoc_sdram_bankmachine5_wrport_dat_w;
wire videosoc_sdram_bankmachine5_do_read;
wire [2:0] videosoc_sdram_bankmachine5_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine5_rdport_dat_r;
wire videosoc_sdram_bankmachine5_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine5_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine5_fifo_in_first;
wire videosoc_sdram_bankmachine5_fifo_in_last;
wire videosoc_sdram_bankmachine5_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine5_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine5_fifo_out_first;
wire videosoc_sdram_bankmachine5_fifo_out_last;
reg videosoc_sdram_bankmachine5_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine5_openrow = 15'd0;
wire videosoc_sdram_bankmachine5_hit;
reg videosoc_sdram_bankmachine5_track_open = 1'd0;
reg videosoc_sdram_bankmachine5_track_close = 1'd0;
reg videosoc_sdram_bankmachine5_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine5_wait;
wire videosoc_sdram_bankmachine5_done;
reg [2:0] videosoc_sdram_bankmachine5_count = 3'd5;
wire videosoc_sdram_bankmachine6_req_valid;
wire videosoc_sdram_bankmachine6_req_ready;
wire videosoc_sdram_bankmachine6_req_we;
wire [21:0] videosoc_sdram_bankmachine6_req_adr;
wire videosoc_sdram_bankmachine6_req_lock;
reg videosoc_sdram_bankmachine6_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine6_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine6_refresh_req;
reg videosoc_sdram_bankmachine6_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine6_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine6_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine6_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine6_cmd_payload_ba;
reg videosoc_sdram_bankmachine6_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine6_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine6_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine6_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine6_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine6_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine6_sink_valid;
wire videosoc_sdram_bankmachine6_sink_ready;
reg videosoc_sdram_bankmachine6_sink_first = 1'd0;
reg videosoc_sdram_bankmachine6_sink_last = 1'd0;
wire videosoc_sdram_bankmachine6_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine6_sink_payload_adr;
wire videosoc_sdram_bankmachine6_source_valid;
wire videosoc_sdram_bankmachine6_source_ready;
wire videosoc_sdram_bankmachine6_source_first;
wire videosoc_sdram_bankmachine6_source_last;
wire videosoc_sdram_bankmachine6_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine6_source_payload_adr;
wire videosoc_sdram_bankmachine6_syncfifo6_we;
wire videosoc_sdram_bankmachine6_syncfifo6_writable;
wire videosoc_sdram_bankmachine6_syncfifo6_re;
wire videosoc_sdram_bankmachine6_syncfifo6_readable;
wire [24:0] videosoc_sdram_bankmachine6_syncfifo6_din;
wire [24:0] videosoc_sdram_bankmachine6_syncfifo6_dout;
reg [3:0] videosoc_sdram_bankmachine6_level = 4'd0;
reg videosoc_sdram_bankmachine6_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine6_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine6_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine6_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine6_wrport_dat_r;
wire videosoc_sdram_bankmachine6_wrport_we;
wire [24:0] videosoc_sdram_bankmachine6_wrport_dat_w;
wire videosoc_sdram_bankmachine6_do_read;
wire [2:0] videosoc_sdram_bankmachine6_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine6_rdport_dat_r;
wire videosoc_sdram_bankmachine6_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine6_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine6_fifo_in_first;
wire videosoc_sdram_bankmachine6_fifo_in_last;
wire videosoc_sdram_bankmachine6_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine6_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine6_fifo_out_first;
wire videosoc_sdram_bankmachine6_fifo_out_last;
reg videosoc_sdram_bankmachine6_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine6_openrow = 15'd0;
wire videosoc_sdram_bankmachine6_hit;
reg videosoc_sdram_bankmachine6_track_open = 1'd0;
reg videosoc_sdram_bankmachine6_track_close = 1'd0;
reg videosoc_sdram_bankmachine6_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine6_wait;
wire videosoc_sdram_bankmachine6_done;
reg [2:0] videosoc_sdram_bankmachine6_count = 3'd5;
wire videosoc_sdram_bankmachine7_req_valid;
wire videosoc_sdram_bankmachine7_req_ready;
wire videosoc_sdram_bankmachine7_req_we;
wire [21:0] videosoc_sdram_bankmachine7_req_adr;
wire videosoc_sdram_bankmachine7_req_lock;
reg videosoc_sdram_bankmachine7_req_wdata_ready = 1'd0;
reg videosoc_sdram_bankmachine7_req_rdata_valid = 1'd0;
wire videosoc_sdram_bankmachine7_refresh_req;
reg videosoc_sdram_bankmachine7_refresh_gnt = 1'd0;
reg videosoc_sdram_bankmachine7_cmd_valid = 1'd0;
reg videosoc_sdram_bankmachine7_cmd_ready = 1'd0;
reg [14:0] videosoc_sdram_bankmachine7_cmd_payload_a = 15'd0;
wire [2:0] videosoc_sdram_bankmachine7_cmd_payload_ba;
reg videosoc_sdram_bankmachine7_cmd_payload_cas = 1'd0;
reg videosoc_sdram_bankmachine7_cmd_payload_ras = 1'd0;
reg videosoc_sdram_bankmachine7_cmd_payload_we = 1'd0;
reg videosoc_sdram_bankmachine7_cmd_payload_is_cmd = 1'd0;
reg videosoc_sdram_bankmachine7_cmd_payload_is_read = 1'd0;
reg videosoc_sdram_bankmachine7_cmd_payload_is_write = 1'd0;
wire videosoc_sdram_bankmachine7_sink_valid;
wire videosoc_sdram_bankmachine7_sink_ready;
reg videosoc_sdram_bankmachine7_sink_first = 1'd0;
reg videosoc_sdram_bankmachine7_sink_last = 1'd0;
wire videosoc_sdram_bankmachine7_sink_payload_we;
wire [21:0] videosoc_sdram_bankmachine7_sink_payload_adr;
wire videosoc_sdram_bankmachine7_source_valid;
wire videosoc_sdram_bankmachine7_source_ready;
wire videosoc_sdram_bankmachine7_source_first;
wire videosoc_sdram_bankmachine7_source_last;
wire videosoc_sdram_bankmachine7_source_payload_we;
wire [21:0] videosoc_sdram_bankmachine7_source_payload_adr;
wire videosoc_sdram_bankmachine7_syncfifo7_we;
wire videosoc_sdram_bankmachine7_syncfifo7_writable;
wire videosoc_sdram_bankmachine7_syncfifo7_re;
wire videosoc_sdram_bankmachine7_syncfifo7_readable;
wire [24:0] videosoc_sdram_bankmachine7_syncfifo7_din;
wire [24:0] videosoc_sdram_bankmachine7_syncfifo7_dout;
reg [3:0] videosoc_sdram_bankmachine7_level = 4'd0;
reg videosoc_sdram_bankmachine7_replace = 1'd0;
reg [2:0] videosoc_sdram_bankmachine7_produce = 3'd0;
reg [2:0] videosoc_sdram_bankmachine7_consume = 3'd0;
reg [2:0] videosoc_sdram_bankmachine7_wrport_adr = 3'd0;
wire [24:0] videosoc_sdram_bankmachine7_wrport_dat_r;
wire videosoc_sdram_bankmachine7_wrport_we;
wire [24:0] videosoc_sdram_bankmachine7_wrport_dat_w;
wire videosoc_sdram_bankmachine7_do_read;
wire [2:0] videosoc_sdram_bankmachine7_rdport_adr;
wire [24:0] videosoc_sdram_bankmachine7_rdport_dat_r;
wire videosoc_sdram_bankmachine7_fifo_in_payload_we;
wire [21:0] videosoc_sdram_bankmachine7_fifo_in_payload_adr;
wire videosoc_sdram_bankmachine7_fifo_in_first;
wire videosoc_sdram_bankmachine7_fifo_in_last;
wire videosoc_sdram_bankmachine7_fifo_out_payload_we;
wire [21:0] videosoc_sdram_bankmachine7_fifo_out_payload_adr;
wire videosoc_sdram_bankmachine7_fifo_out_first;
wire videosoc_sdram_bankmachine7_fifo_out_last;
reg videosoc_sdram_bankmachine7_has_openrow = 1'd0;
reg [14:0] videosoc_sdram_bankmachine7_openrow = 15'd0;
wire videosoc_sdram_bankmachine7_hit;
reg videosoc_sdram_bankmachine7_track_open = 1'd0;
reg videosoc_sdram_bankmachine7_track_close = 1'd0;
reg videosoc_sdram_bankmachine7_sel_row_adr = 1'd0;
wire videosoc_sdram_bankmachine7_wait;
wire videosoc_sdram_bankmachine7_done;
reg [2:0] videosoc_sdram_bankmachine7_count = 3'd5;
reg videosoc_sdram_choose_cmd_want_reads = 1'd0;
reg videosoc_sdram_choose_cmd_want_writes = 1'd0;
reg videosoc_sdram_choose_cmd_want_cmds = 1'd0;
wire videosoc_sdram_choose_cmd_cmd_valid;
reg videosoc_sdram_choose_cmd_cmd_ready = 1'd0;
wire [14:0] videosoc_sdram_choose_cmd_cmd_payload_a;
wire [2:0] videosoc_sdram_choose_cmd_cmd_payload_ba;
reg videosoc_sdram_choose_cmd_cmd_payload_cas = 1'd0;
reg videosoc_sdram_choose_cmd_cmd_payload_ras = 1'd0;
reg videosoc_sdram_choose_cmd_cmd_payload_we = 1'd0;
wire videosoc_sdram_choose_cmd_cmd_payload_is_cmd;
wire videosoc_sdram_choose_cmd_cmd_payload_is_read;
wire videosoc_sdram_choose_cmd_cmd_payload_is_write;
reg [7:0] videosoc_sdram_choose_cmd_valids = 8'd0;
wire [7:0] videosoc_sdram_choose_cmd_request;
reg [2:0] videosoc_sdram_choose_cmd_grant = 3'd0;
wire videosoc_sdram_choose_cmd_ce;
reg videosoc_sdram_choose_req_want_reads = 1'd0;
reg videosoc_sdram_choose_req_want_writes = 1'd0;
reg videosoc_sdram_choose_req_want_cmds = 1'd0;
wire videosoc_sdram_choose_req_cmd_valid;
reg videosoc_sdram_choose_req_cmd_ready = 1'd0;
wire [14:0] videosoc_sdram_choose_req_cmd_payload_a;
wire [2:0] videosoc_sdram_choose_req_cmd_payload_ba;
reg videosoc_sdram_choose_req_cmd_payload_cas = 1'd0;
reg videosoc_sdram_choose_req_cmd_payload_ras = 1'd0;
reg videosoc_sdram_choose_req_cmd_payload_we = 1'd0;
wire videosoc_sdram_choose_req_cmd_payload_is_cmd;
wire videosoc_sdram_choose_req_cmd_payload_is_read;
wire videosoc_sdram_choose_req_cmd_payload_is_write;
reg [7:0] videosoc_sdram_choose_req_valids = 8'd0;
wire [7:0] videosoc_sdram_choose_req_request;
reg [2:0] videosoc_sdram_choose_req_grant = 3'd0;
wire videosoc_sdram_choose_req_ce;
reg [14:0] videosoc_sdram_nop_a = 15'd0;
reg [2:0] videosoc_sdram_nop_ba = 3'd0;
reg videosoc_sdram_nop_cas = 1'd0;
reg videosoc_sdram_nop_ras = 1'd0;
reg videosoc_sdram_nop_we = 1'd0;
reg [1:0] videosoc_sdram_sel0 = 2'd0;
reg [1:0] videosoc_sdram_sel1 = 2'd0;
reg [1:0] videosoc_sdram_sel2 = 2'd0;
reg [1:0] videosoc_sdram_sel3 = 2'd0;
wire videosoc_sdram_read_available;
wire videosoc_sdram_write_available;
reg videosoc_sdram_en0 = 1'd0;
wire videosoc_sdram_max_time0;
reg [4:0] videosoc_sdram_time0 = 5'd0;
reg videosoc_sdram_en1 = 1'd0;
wire videosoc_sdram_max_time1;
reg [3:0] videosoc_sdram_time1 = 4'd0;
wire videosoc_sdram_go_to_refresh;
wire videosoc_sdram_bandwidth_update_re;
wire videosoc_sdram_bandwidth_update_r;
reg videosoc_sdram_bandwidth_update_w = 1'd0;
reg [23:0] videosoc_sdram_bandwidth_nreads_status = 24'd0;
reg [23:0] videosoc_sdram_bandwidth_nwrites_status = 24'd0;
reg [7:0] videosoc_sdram_bandwidth_data_width_status = 8'd128;
reg videosoc_sdram_bandwidth_cmd_valid = 1'd0;
reg videosoc_sdram_bandwidth_cmd_ready = 1'd0;
reg videosoc_sdram_bandwidth_cmd_is_read = 1'd0;
reg videosoc_sdram_bandwidth_cmd_is_write = 1'd0;
reg [23:0] videosoc_sdram_bandwidth_counter = 24'd0;
reg videosoc_sdram_bandwidth_period = 1'd0;
reg [23:0] videosoc_sdram_bandwidth_nreads = 24'd0;
reg [23:0] videosoc_sdram_bandwidth_nwrites = 24'd0;
reg [23:0] videosoc_sdram_bandwidth_nreads_r = 24'd0;
reg [23:0] videosoc_sdram_bandwidth_nwrites_r = 24'd0;
wire [29:0] videosoc_interface1_wb_sdram_adr;
wire [31:0] videosoc_interface1_wb_sdram_dat_w;
wire [31:0] videosoc_interface1_wb_sdram_dat_r;
wire [3:0] videosoc_interface1_wb_sdram_sel;
wire videosoc_interface1_wb_sdram_cyc;
wire videosoc_interface1_wb_sdram_stb;
wire videosoc_interface1_wb_sdram_ack;
wire videosoc_interface1_wb_sdram_we;
wire [2:0] videosoc_interface1_wb_sdram_cti;
wire [1:0] videosoc_interface1_wb_sdram_bte;
wire videosoc_interface1_wb_sdram_err;
reg videosoc_port_cmd_valid = 1'd0;
wire videosoc_port_cmd_ready;
reg videosoc_port_cmd_payload_we = 1'd0;
wire [24:0] videosoc_port_cmd_payload_adr;
reg videosoc_port_wdata_valid = 1'd0;
wire videosoc_port_wdata_ready;
wire [127:0] videosoc_port_wdata_payload_data;
wire [15:0] videosoc_port_wdata_payload_we;
wire videosoc_port_rdata_valid;
reg videosoc_port_rdata_ready = 1'd0;
wire [127:0] videosoc_port_rdata_payload_data;
wire [29:0] videosoc_interface_adr;
wire [127:0] videosoc_interface_dat_w;
wire [127:0] videosoc_interface_dat_r;
wire [15:0] videosoc_interface_sel;
reg videosoc_interface_cyc = 1'd0;
reg videosoc_interface_stb = 1'd0;
reg videosoc_interface_ack = 1'd0;
reg videosoc_interface_we = 1'd0;
wire [8:0] videosoc_data_port_adr;
wire [127:0] videosoc_data_port_dat_r;
reg [15:0] videosoc_data_port_we = 16'd0;
reg [127:0] videosoc_data_port_dat_w = 128'd0;
reg videosoc_write_from_slave = 1'd0;
reg [1:0] videosoc_adr_offset_r = 2'd0;
wire [8:0] videosoc_tag_port_adr;
wire [23:0] videosoc_tag_port_dat_r;
reg videosoc_tag_port_we = 1'd0;
wire [23:0] videosoc_tag_port_dat_w;
wire [22:0] videosoc_tag_do_tag;
wire videosoc_tag_do_dirty;
wire [22:0] videosoc_tag_di_tag;
reg videosoc_tag_di_dirty = 1'd0;
reg videosoc_word_clr = 1'd0;
reg videosoc_word_inc = 1'd0;
reg videosoc_clk0 = 1'd0;
wire [29:0] videosoc_bus_adr;
wire [31:0] videosoc_bus_dat_w;
wire [31:0] videosoc_bus_dat_r;
wire [3:0] videosoc_bus_sel;
wire videosoc_bus_cyc;
wire videosoc_bus_stb;
reg videosoc_bus_ack = 1'd0;
wire videosoc_bus_we;
wire [2:0] videosoc_bus_cti;
wire [1:0] videosoc_bus_bte;
reg videosoc_bus_err = 1'd0;
reg [3:0] videosoc_bitbang_storage_full = 4'd0;
wire [3:0] videosoc_bitbang_storage;
reg videosoc_bitbang_re = 1'd0;
reg videosoc_miso_status = 1'd0;
reg videosoc_bitbang_en_storage_full = 1'd0;
wire videosoc_bitbang_en_storage;
reg videosoc_bitbang_en_re = 1'd0;
reg videosoc_cs_n = 1'd1;
reg videosoc_clk1 = 1'd0;
reg [31:0] videosoc_sr = 32'd0;
reg videosoc_i = 1'd0;
reg videosoc_miso = 1'd0;
reg [7:0] videosoc_counter = 8'd0;
reg ethphy_reset_storage_full = 1'd0;
wire ethphy_reset_storage;
reg ethphy_reset_re = 1'd0;
(* dont_touch = "true" *) wire eth_rx_clk;
wire eth_rx_rst;
(* dont_touch = "true" *) wire eth_tx_clk;
wire eth_tx_rst;
wire eth_tx90_clk;
wire ethphy_eth_rx_clk_ibuf;
wire ethphy_pll_locked;
wire ethphy_pll_fb;
wire ethphy_pll_clk_tx;
wire ethphy_pll_clk_tx90;
wire ethphy_eth_tx_clk_obuf;
(* ars_false_path = "true" *) wire ethphy_reset0;
wire ethphy_reset1;
reg [8:0] ethphy_counter = 9'd0;
wire ethphy_counter_done;
wire ethphy_counter_ce;
wire ethphy_sink_valid;
wire ethphy_sink_ready;
wire ethphy_sink_first;
wire ethphy_sink_last;
wire [7:0] ethphy_sink_payload_data;
wire ethphy_sink_payload_last_be;
wire ethphy_sink_payload_error;
wire ethphy_tx_ctl_obuf;
wire [3:0] ethphy_tx_data_obuf;
reg ethphy_source_valid = 1'd0;
wire ethphy_source_ready;
reg ethphy_source_first = 1'd0;
wire ethphy_source_last;
reg [7:0] ethphy_source_payload_data = 8'd0;
reg ethphy_source_payload_last_be = 1'd0;
reg ethphy_source_payload_error = 1'd0;
wire ethphy_rx_ctl_ibuf;
wire ethphy_rx_ctl_idelay;
wire ethphy_rx_ctl;
wire [3:0] ethphy_rx_data_ibuf;
wire [3:0] ethphy_rx_data_idelay;
wire [7:0] ethphy_rx_data;
reg ethphy_rx_ctl_d = 1'd0;
wire ethphy_last;
reg [2:0] ethphy_storage_full = 3'd0;
wire [2:0] ethphy_storage;
reg ethphy_re = 1'd0;
wire ethphy_status;
wire ethphy_data_w;
wire ethphy_data_oe;
wire ethphy_data_r;
wire ethmac_tx_gap_inserter_sink_valid;
reg ethmac_tx_gap_inserter_sink_ready = 1'd0;
wire ethmac_tx_gap_inserter_sink_first;
wire ethmac_tx_gap_inserter_sink_last;
wire [7:0] ethmac_tx_gap_inserter_sink_payload_data;
wire ethmac_tx_gap_inserter_sink_payload_last_be;
wire ethmac_tx_gap_inserter_sink_payload_error;
reg ethmac_tx_gap_inserter_source_valid = 1'd0;
wire ethmac_tx_gap_inserter_source_ready;
reg ethmac_tx_gap_inserter_source_first = 1'd0;
reg ethmac_tx_gap_inserter_source_last = 1'd0;
reg [7:0] ethmac_tx_gap_inserter_source_payload_data = 8'd0;
reg ethmac_tx_gap_inserter_source_payload_last_be = 1'd0;
reg ethmac_tx_gap_inserter_source_payload_error = 1'd0;
reg [3:0] ethmac_tx_gap_inserter_counter = 4'd0;
reg ethmac_tx_gap_inserter_counter_reset = 1'd0;
reg ethmac_tx_gap_inserter_counter_ce = 1'd0;
reg ethmac_preamble_crc_status = 1'd1;
reg [31:0] ethmac_preamble_errors_status = 32'd0;
reg [31:0] ethmac_crc_errors_status = 32'd0;
wire ethmac_preamble_inserter_sink_valid;
reg ethmac_preamble_inserter_sink_ready = 1'd0;
wire ethmac_preamble_inserter_sink_first;
wire ethmac_preamble_inserter_sink_last;
wire [7:0] ethmac_preamble_inserter_sink_payload_data;
wire ethmac_preamble_inserter_sink_payload_last_be;
wire ethmac_preamble_inserter_sink_payload_error;
reg ethmac_preamble_inserter_source_valid = 1'd0;
wire ethmac_preamble_inserter_source_ready;
reg ethmac_preamble_inserter_source_first = 1'd0;
reg ethmac_preamble_inserter_source_last = 1'd0;
reg [7:0] ethmac_preamble_inserter_source_payload_data = 8'd0;
wire ethmac_preamble_inserter_source_payload_last_be;
reg ethmac_preamble_inserter_source_payload_error = 1'd0;
reg [63:0] ethmac_preamble_inserter_preamble = 64'd15372286728091293013;
reg [2:0] ethmac_preamble_inserter_cnt = 3'd0;
reg ethmac_preamble_inserter_clr_cnt = 1'd0;
reg ethmac_preamble_inserter_inc_cnt = 1'd0;
wire ethmac_preamble_checker_sink_valid;
reg ethmac_preamble_checker_sink_ready = 1'd0;
wire ethmac_preamble_checker_sink_first;
wire ethmac_preamble_checker_sink_last;
wire [7:0] ethmac_preamble_checker_sink_payload_data;
wire ethmac_preamble_checker_sink_payload_last_be;
wire ethmac_preamble_checker_sink_payload_error;
reg ethmac_preamble_checker_source_valid = 1'd0;
wire ethmac_preamble_checker_source_ready;
reg ethmac_preamble_checker_source_first = 1'd0;
reg ethmac_preamble_checker_source_last = 1'd0;
wire [7:0] ethmac_preamble_checker_source_payload_data;
wire ethmac_preamble_checker_source_payload_last_be;
reg ethmac_preamble_checker_source_payload_error = 1'd0;
reg ethmac_preamble_checker_error = 1'd0;
wire ethmac_crc32_inserter_sink_valid;
reg ethmac_crc32_inserter_sink_ready = 1'd0;
wire ethmac_crc32_inserter_sink_first;
wire ethmac_crc32_inserter_sink_last;
wire [7:0] ethmac_crc32_inserter_sink_payload_data;
wire ethmac_crc32_inserter_sink_payload_last_be;
wire ethmac_crc32_inserter_sink_payload_error;
reg ethmac_crc32_inserter_source_valid = 1'd0;
wire ethmac_crc32_inserter_source_ready;
reg ethmac_crc32_inserter_source_first = 1'd0;
reg ethmac_crc32_inserter_source_last = 1'd0;
reg [7:0] ethmac_crc32_inserter_source_payload_data = 8'd0;
reg ethmac_crc32_inserter_source_payload_last_be = 1'd0;
reg ethmac_crc32_inserter_source_payload_error = 1'd0;
reg [7:0] ethmac_crc32_inserter_data0 = 8'd0;
wire [31:0] ethmac_crc32_inserter_value;
wire ethmac_crc32_inserter_error;
wire [7:0] ethmac_crc32_inserter_data1;
wire [31:0] ethmac_crc32_inserter_last;
reg [31:0] ethmac_crc32_inserter_next = 32'd0;
reg [31:0] ethmac_crc32_inserter_reg = 32'd4294967295;
reg ethmac_crc32_inserter_ce = 1'd0;
reg ethmac_crc32_inserter_reset = 1'd0;
reg [1:0] ethmac_crc32_inserter_cnt = 2'd3;
wire ethmac_crc32_inserter_cnt_done;
reg ethmac_crc32_inserter_is_ongoing0 = 1'd0;
reg ethmac_crc32_inserter_is_ongoing1 = 1'd0;
wire ethmac_crc32_checker_sink_sink_valid;
reg ethmac_crc32_checker_sink_sink_ready = 1'd0;
wire ethmac_crc32_checker_sink_sink_first;
wire ethmac_crc32_checker_sink_sink_last;
wire [7:0] ethmac_crc32_checker_sink_sink_payload_data;
wire ethmac_crc32_checker_sink_sink_payload_last_be;
wire ethmac_crc32_checker_sink_sink_payload_error;
wire ethmac_crc32_checker_source_source_valid;
wire ethmac_crc32_checker_source_source_ready;
reg ethmac_crc32_checker_source_source_first = 1'd0;
wire ethmac_crc32_checker_source_source_last;
wire [7:0] ethmac_crc32_checker_source_source_payload_data;
wire ethmac_crc32_checker_source_source_payload_last_be;
reg ethmac_crc32_checker_source_source_payload_error = 1'd0;
wire ethmac_crc32_checker_error;
wire [7:0] ethmac_crc32_checker_crc_data0;
wire [31:0] ethmac_crc32_checker_crc_value;
wire ethmac_crc32_checker_crc_error;
wire [7:0] ethmac_crc32_checker_crc_data1;
wire [31:0] ethmac_crc32_checker_crc_last;
reg [31:0] ethmac_crc32_checker_crc_next = 32'd0;
reg [31:0] ethmac_crc32_checker_crc_reg = 32'd4294967295;
reg ethmac_crc32_checker_crc_ce = 1'd0;
reg ethmac_crc32_checker_crc_reset = 1'd0;
reg ethmac_crc32_checker_syncfifo_sink_valid = 1'd0;
wire ethmac_crc32_checker_syncfifo_sink_ready;
wire ethmac_crc32_checker_syncfifo_sink_first;
wire ethmac_crc32_checker_syncfifo_sink_last;
wire [7:0] ethmac_crc32_checker_syncfifo_sink_payload_data;
wire ethmac_crc32_checker_syncfifo_sink_payload_last_be;
wire ethmac_crc32_checker_syncfifo_sink_payload_error;
wire ethmac_crc32_checker_syncfifo_source_valid;
wire ethmac_crc32_checker_syncfifo_source_ready;
wire ethmac_crc32_checker_syncfifo_source_first;
wire ethmac_crc32_checker_syncfifo_source_last;
wire [7:0] ethmac_crc32_checker_syncfifo_source_payload_data;
wire ethmac_crc32_checker_syncfifo_source_payload_last_be;
wire ethmac_crc32_checker_syncfifo_source_payload_error;
wire ethmac_crc32_checker_syncfifo_syncfifo_we;
wire ethmac_crc32_checker_syncfifo_syncfifo_writable;
wire ethmac_crc32_checker_syncfifo_syncfifo_re;
wire ethmac_crc32_checker_syncfifo_syncfifo_readable;
wire [11:0] ethmac_crc32_checker_syncfifo_syncfifo_din;
wire [11:0] ethmac_crc32_checker_syncfifo_syncfifo_dout;
reg [2:0] ethmac_crc32_checker_syncfifo_level = 3'd0;
reg ethmac_crc32_checker_syncfifo_replace = 1'd0;
reg [2:0] ethmac_crc32_checker_syncfifo_produce = 3'd0;
reg [2:0] ethmac_crc32_checker_syncfifo_consume = 3'd0;
reg [2:0] ethmac_crc32_checker_syncfifo_wrport_adr = 3'd0;
wire [11:0] ethmac_crc32_checker_syncfifo_wrport_dat_r;
wire ethmac_crc32_checker_syncfifo_wrport_we;
wire [11:0] ethmac_crc32_checker_syncfifo_wrport_dat_w;
wire ethmac_crc32_checker_syncfifo_do_read;
wire [2:0] ethmac_crc32_checker_syncfifo_rdport_adr;
wire [11:0] ethmac_crc32_checker_syncfifo_rdport_dat_r;
wire [7:0] ethmac_crc32_checker_syncfifo_fifo_in_payload_data;
wire ethmac_crc32_checker_syncfifo_fifo_in_payload_last_be;
wire ethmac_crc32_checker_syncfifo_fifo_in_payload_error;
wire ethmac_crc32_checker_syncfifo_fifo_in_first;
wire ethmac_crc32_checker_syncfifo_fifo_in_last;
wire [7:0] ethmac_crc32_checker_syncfifo_fifo_out_payload_data;
wire ethmac_crc32_checker_syncfifo_fifo_out_payload_last_be;
wire ethmac_crc32_checker_syncfifo_fifo_out_payload_error;
wire ethmac_crc32_checker_syncfifo_fifo_out_first;
wire ethmac_crc32_checker_syncfifo_fifo_out_last;
reg ethmac_crc32_checker_fifo_reset = 1'd0;
wire ethmac_crc32_checker_fifo_in;
wire ethmac_crc32_checker_fifo_out;
wire ethmac_crc32_checker_fifo_full;
wire ethmac_ps_preamble_error_i;
wire ethmac_ps_preamble_error_o;
reg ethmac_ps_preamble_error_toggle_i = 1'd0;
wire ethmac_ps_preamble_error_toggle_o;
reg ethmac_ps_preamble_error_toggle_o_r = 1'd0;
wire ethmac_ps_crc_error_i;
wire ethmac_ps_crc_error_o;
reg ethmac_ps_crc_error_toggle_i = 1'd0;
wire ethmac_ps_crc_error_toggle_o;
reg ethmac_ps_crc_error_toggle_o_r = 1'd0;
wire ethmac_padding_inserter_sink_valid;
reg ethmac_padding_inserter_sink_ready = 1'd0;
wire ethmac_padding_inserter_sink_first;
wire ethmac_padding_inserter_sink_last;
wire [7:0] ethmac_padding_inserter_sink_payload_data;
wire ethmac_padding_inserter_sink_payload_last_be;
wire ethmac_padding_inserter_sink_payload_error;
reg ethmac_padding_inserter_source_valid = 1'd0;
wire ethmac_padding_inserter_source_ready;
reg ethmac_padding_inserter_source_first = 1'd0;
reg ethmac_padding_inserter_source_last = 1'd0;
reg [7:0] ethmac_padding_inserter_source_payload_data = 8'd0;
reg ethmac_padding_inserter_source_payload_last_be = 1'd0;
reg ethmac_padding_inserter_source_payload_error = 1'd0;
reg [15:0] ethmac_padding_inserter_counter = 16'd1;
wire ethmac_padding_inserter_counter_done;
reg ethmac_padding_inserter_counter_reset = 1'd0;
reg ethmac_padding_inserter_counter_ce = 1'd0;
wire ethmac_padding_checker_sink_valid;
wire ethmac_padding_checker_sink_ready;
wire ethmac_padding_checker_sink_first;
wire ethmac_padding_checker_sink_last;
wire [7:0] ethmac_padding_checker_sink_payload_data;
wire ethmac_padding_checker_sink_payload_last_be;
wire ethmac_padding_checker_sink_payload_error;
wire ethmac_padding_checker_source_valid;
wire ethmac_padding_checker_source_ready;
wire ethmac_padding_checker_source_first;
wire ethmac_padding_checker_source_last;
wire [7:0] ethmac_padding_checker_source_payload_data;
wire ethmac_padding_checker_source_payload_last_be;
wire ethmac_padding_checker_source_payload_error;
wire ethmac_tx_last_be_sink_valid;
wire ethmac_tx_last_be_sink_ready;
wire ethmac_tx_last_be_sink_first;
wire ethmac_tx_last_be_sink_last;
wire [7:0] ethmac_tx_last_be_sink_payload_data;
wire ethmac_tx_last_be_sink_payload_last_be;
wire ethmac_tx_last_be_sink_payload_error;
wire ethmac_tx_last_be_source_valid;
wire ethmac_tx_last_be_source_ready;
reg ethmac_tx_last_be_source_first = 1'd0;
wire ethmac_tx_last_be_source_last;
wire [7:0] ethmac_tx_last_be_source_payload_data;
reg ethmac_tx_last_be_source_payload_last_be = 1'd0;
reg ethmac_tx_last_be_source_payload_error = 1'd0;
reg ethmac_tx_last_be_ongoing = 1'd1;
wire ethmac_rx_last_be_sink_valid;
wire ethmac_rx_last_be_sink_ready;
wire ethmac_rx_last_be_sink_first;
wire ethmac_rx_last_be_sink_last;
wire [7:0] ethmac_rx_last_be_sink_payload_data;
wire ethmac_rx_last_be_sink_payload_last_be;
wire ethmac_rx_last_be_sink_payload_error;
wire ethmac_rx_last_be_source_valid;
wire ethmac_rx_last_be_source_ready;
wire ethmac_rx_last_be_source_first;
wire ethmac_rx_last_be_source_last;
wire [7:0] ethmac_rx_last_be_source_payload_data;
reg ethmac_rx_last_be_source_payload_last_be = 1'd0;
wire ethmac_rx_last_be_source_payload_error;
wire ethmac_tx_converter_sink_valid;
wire ethmac_tx_converter_sink_ready;
wire ethmac_tx_converter_sink_first;
wire ethmac_tx_converter_sink_last;
wire [31:0] ethmac_tx_converter_sink_payload_data;
wire [3:0] ethmac_tx_converter_sink_payload_last_be;
wire [3:0] ethmac_tx_converter_sink_payload_error;
wire ethmac_tx_converter_source_valid;
wire ethmac_tx_converter_source_ready;
wire ethmac_tx_converter_source_first;
wire ethmac_tx_converter_source_last;
wire [7:0] ethmac_tx_converter_source_payload_data;
wire ethmac_tx_converter_source_payload_last_be;
wire ethmac_tx_converter_source_payload_error;
wire ethmac_tx_converter_converter_sink_valid;
wire ethmac_tx_converter_converter_sink_ready;
wire ethmac_tx_converter_converter_sink_first;
wire ethmac_tx_converter_converter_sink_last;
reg [39:0] ethmac_tx_converter_converter_sink_payload_data = 40'd0;
wire ethmac_tx_converter_converter_source_valid;
wire ethmac_tx_converter_converter_source_ready;
wire ethmac_tx_converter_converter_source_first;
wire ethmac_tx_converter_converter_source_last;
reg [9:0] ethmac_tx_converter_converter_source_payload_data = 10'd0;
wire ethmac_tx_converter_converter_source_payload_valid_token_count;
reg [1:0] ethmac_tx_converter_converter_mux = 2'd0;
wire ethmac_tx_converter_converter_first;
wire ethmac_tx_converter_converter_last;
wire ethmac_tx_converter_source_source_valid;
wire ethmac_tx_converter_source_source_ready;
wire ethmac_tx_converter_source_source_first;
wire ethmac_tx_converter_source_source_last;
wire [9:0] ethmac_tx_converter_source_source_payload_data;
wire ethmac_rx_converter_sink_valid;
wire ethmac_rx_converter_sink_ready;
wire ethmac_rx_converter_sink_first;
wire ethmac_rx_converter_sink_last;
wire [7:0] ethmac_rx_converter_sink_payload_data;
wire ethmac_rx_converter_sink_payload_last_be;
wire ethmac_rx_converter_sink_payload_error;
wire ethmac_rx_converter_source_valid;
wire ethmac_rx_converter_source_ready;
wire ethmac_rx_converter_source_first;
wire ethmac_rx_converter_source_last;
reg [31:0] ethmac_rx_converter_source_payload_data = 32'd0;
reg [3:0] ethmac_rx_converter_source_payload_last_be = 4'd0;
reg [3:0] ethmac_rx_converter_source_payload_error = 4'd0;
wire ethmac_rx_converter_converter_sink_valid;
wire ethmac_rx_converter_converter_sink_ready;
wire ethmac_rx_converter_converter_sink_first;
wire ethmac_rx_converter_converter_sink_last;
wire [9:0] ethmac_rx_converter_converter_sink_payload_data;
wire ethmac_rx_converter_converter_source_valid;
wire ethmac_rx_converter_converter_source_ready;
reg ethmac_rx_converter_converter_source_first = 1'd0;
reg ethmac_rx_converter_converter_source_last = 1'd0;
reg [39:0] ethmac_rx_converter_converter_source_payload_data = 40'd0;
reg [2:0] ethmac_rx_converter_converter_source_payload_valid_token_count = 3'd0;
reg [1:0] ethmac_rx_converter_converter_demux = 2'd0;
wire ethmac_rx_converter_converter_load_part;
reg ethmac_rx_converter_converter_strobe_all = 1'd0;
wire ethmac_rx_converter_source_source_valid;
wire ethmac_rx_converter_source_source_ready;
wire ethmac_rx_converter_source_source_first;
wire ethmac_rx_converter_source_source_last;
wire [39:0] ethmac_rx_converter_source_source_payload_data;
wire ethmac_tx_cdc_sink_valid;
wire ethmac_tx_cdc_sink_ready;
wire ethmac_tx_cdc_sink_first;
wire ethmac_tx_cdc_sink_last;
wire [31:0] ethmac_tx_cdc_sink_payload_data;
wire [3:0] ethmac_tx_cdc_sink_payload_last_be;
wire [3:0] ethmac_tx_cdc_sink_payload_error;
wire ethmac_tx_cdc_source_valid;
wire ethmac_tx_cdc_source_ready;
wire ethmac_tx_cdc_source_first;
wire ethmac_tx_cdc_source_last;
wire [31:0] ethmac_tx_cdc_source_payload_data;
wire [3:0] ethmac_tx_cdc_source_payload_last_be;
wire [3:0] ethmac_tx_cdc_source_payload_error;
wire ethmac_tx_cdc_asyncfifo_we;
wire ethmac_tx_cdc_asyncfifo_writable;
wire ethmac_tx_cdc_asyncfifo_re;
wire ethmac_tx_cdc_asyncfifo_readable;
wire [41:0] ethmac_tx_cdc_asyncfifo_din;
wire [41:0] ethmac_tx_cdc_asyncfifo_dout;
wire ethmac_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] ethmac_tx_cdc_graycounter0_q = 7'd0;
wire [6:0] ethmac_tx_cdc_graycounter0_q_next;
reg [6:0] ethmac_tx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] ethmac_tx_cdc_graycounter0_q_next_binary = 7'd0;
wire ethmac_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] ethmac_tx_cdc_graycounter1_q = 7'd0;
wire [6:0] ethmac_tx_cdc_graycounter1_q_next;
reg [6:0] ethmac_tx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] ethmac_tx_cdc_graycounter1_q_next_binary = 7'd0;
wire [6:0] ethmac_tx_cdc_produce_rdomain;
wire [6:0] ethmac_tx_cdc_consume_wdomain;
wire [5:0] ethmac_tx_cdc_wrport_adr;
wire [41:0] ethmac_tx_cdc_wrport_dat_r;
wire ethmac_tx_cdc_wrport_we;
wire [41:0] ethmac_tx_cdc_wrport_dat_w;
wire [5:0] ethmac_tx_cdc_rdport_adr;
wire [41:0] ethmac_tx_cdc_rdport_dat_r;
wire [31:0] ethmac_tx_cdc_fifo_in_payload_data;
wire [3:0] ethmac_tx_cdc_fifo_in_payload_last_be;
wire [3:0] ethmac_tx_cdc_fifo_in_payload_error;
wire ethmac_tx_cdc_fifo_in_first;
wire ethmac_tx_cdc_fifo_in_last;
wire [31:0] ethmac_tx_cdc_fifo_out_payload_data;
wire [3:0] ethmac_tx_cdc_fifo_out_payload_last_be;
wire [3:0] ethmac_tx_cdc_fifo_out_payload_error;
wire ethmac_tx_cdc_fifo_out_first;
wire ethmac_tx_cdc_fifo_out_last;
wire ethmac_rx_cdc_sink_valid;
wire ethmac_rx_cdc_sink_ready;
wire ethmac_rx_cdc_sink_first;
wire ethmac_rx_cdc_sink_last;
wire [31:0] ethmac_rx_cdc_sink_payload_data;
wire [3:0] ethmac_rx_cdc_sink_payload_last_be;
wire [3:0] ethmac_rx_cdc_sink_payload_error;
wire ethmac_rx_cdc_source_valid;
wire ethmac_rx_cdc_source_ready;
wire ethmac_rx_cdc_source_first;
wire ethmac_rx_cdc_source_last;
wire [31:0] ethmac_rx_cdc_source_payload_data;
wire [3:0] ethmac_rx_cdc_source_payload_last_be;
wire [3:0] ethmac_rx_cdc_source_payload_error;
wire ethmac_rx_cdc_asyncfifo_we;
wire ethmac_rx_cdc_asyncfifo_writable;
wire ethmac_rx_cdc_asyncfifo_re;
wire ethmac_rx_cdc_asyncfifo_readable;
wire [41:0] ethmac_rx_cdc_asyncfifo_din;
wire [41:0] ethmac_rx_cdc_asyncfifo_dout;
wire ethmac_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] ethmac_rx_cdc_graycounter0_q = 7'd0;
wire [6:0] ethmac_rx_cdc_graycounter0_q_next;
reg [6:0] ethmac_rx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] ethmac_rx_cdc_graycounter0_q_next_binary = 7'd0;
wire ethmac_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] ethmac_rx_cdc_graycounter1_q = 7'd0;
wire [6:0] ethmac_rx_cdc_graycounter1_q_next;
reg [6:0] ethmac_rx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] ethmac_rx_cdc_graycounter1_q_next_binary = 7'd0;
wire [6:0] ethmac_rx_cdc_produce_rdomain;
wire [6:0] ethmac_rx_cdc_consume_wdomain;
wire [5:0] ethmac_rx_cdc_wrport_adr;
wire [41:0] ethmac_rx_cdc_wrport_dat_r;
wire ethmac_rx_cdc_wrport_we;
wire [41:0] ethmac_rx_cdc_wrport_dat_w;
wire [5:0] ethmac_rx_cdc_rdport_adr;
wire [41:0] ethmac_rx_cdc_rdport_dat_r;
wire [31:0] ethmac_rx_cdc_fifo_in_payload_data;
wire [3:0] ethmac_rx_cdc_fifo_in_payload_last_be;
wire [3:0] ethmac_rx_cdc_fifo_in_payload_error;
wire ethmac_rx_cdc_fifo_in_first;
wire ethmac_rx_cdc_fifo_in_last;
wire [31:0] ethmac_rx_cdc_fifo_out_payload_data;
wire [3:0] ethmac_rx_cdc_fifo_out_payload_last_be;
wire [3:0] ethmac_rx_cdc_fifo_out_payload_error;
wire ethmac_rx_cdc_fifo_out_first;
wire ethmac_rx_cdc_fifo_out_last;
wire ethmac_sink_valid;
wire ethmac_sink_ready;
wire ethmac_sink_first;
wire ethmac_sink_last;
wire [31:0] ethmac_sink_payload_data;
wire [3:0] ethmac_sink_payload_last_be;
wire [3:0] ethmac_sink_payload_error;
wire ethmac_source_valid;
wire ethmac_source_ready;
wire ethmac_source_first;
wire ethmac_source_last;
wire [31:0] ethmac_source_payload_data;
wire [3:0] ethmac_source_payload_last_be;
wire [3:0] ethmac_source_payload_error;
wire [29:0] ethmac_bus_adr;
wire [31:0] ethmac_bus_dat_w;
wire [31:0] ethmac_bus_dat_r;
wire [3:0] ethmac_bus_sel;
wire ethmac_bus_cyc;
wire ethmac_bus_stb;
wire ethmac_bus_ack;
wire ethmac_bus_we;
wire [2:0] ethmac_bus_cti;
wire [1:0] ethmac_bus_bte;
wire ethmac_bus_err;
wire ethmac_writer_sink_sink_valid;
reg ethmac_writer_sink_sink_ready = 1'd1;
wire ethmac_writer_sink_sink_first;
wire ethmac_writer_sink_sink_last;
wire [31:0] ethmac_writer_sink_sink_payload_data;
wire [3:0] ethmac_writer_sink_sink_payload_last_be;
wire [3:0] ethmac_writer_sink_sink_payload_error;
wire ethmac_writer_slot_status;
wire [31:0] ethmac_writer_length_status;
reg [31:0] ethmac_writer_errors_status = 32'd0;
wire ethmac_writer_irq;
wire ethmac_writer_available_status;
wire ethmac_writer_available_pending;
wire ethmac_writer_available_trigger;
reg ethmac_writer_available_clear = 1'd0;
wire ethmac_writer_status_re;
wire ethmac_writer_status_r;
wire ethmac_writer_status_w;
wire ethmac_writer_pending_re;
wire ethmac_writer_pending_r;
wire ethmac_writer_pending_w;
reg ethmac_writer_storage_full = 1'd0;
wire ethmac_writer_storage;
reg ethmac_writer_re = 1'd0;
reg [2:0] ethmac_writer_increment = 3'd0;
reg [31:0] ethmac_writer_counter = 32'd0;
reg ethmac_writer_counter_reset = 1'd0;
reg ethmac_writer_counter_ce = 1'd0;
reg ethmac_writer_slot = 1'd0;
reg ethmac_writer_slot_ce = 1'd0;
reg ethmac_writer_ongoing = 1'd0;
reg ethmac_writer_fifo_sink_valid = 1'd0;
wire ethmac_writer_fifo_sink_ready;
reg ethmac_writer_fifo_sink_first = 1'd0;
reg ethmac_writer_fifo_sink_last = 1'd0;
wire ethmac_writer_fifo_sink_payload_slot;
wire [31:0] ethmac_writer_fifo_sink_payload_length;
wire ethmac_writer_fifo_source_valid;
wire ethmac_writer_fifo_source_ready;
wire ethmac_writer_fifo_source_first;
wire ethmac_writer_fifo_source_last;
wire ethmac_writer_fifo_source_payload_slot;
wire [31:0] ethmac_writer_fifo_source_payload_length;
wire ethmac_writer_fifo_syncfifo_we;
wire ethmac_writer_fifo_syncfifo_writable;
wire ethmac_writer_fifo_syncfifo_re;
wire ethmac_writer_fifo_syncfifo_readable;
wire [34:0] ethmac_writer_fifo_syncfifo_din;
wire [34:0] ethmac_writer_fifo_syncfifo_dout;
reg [1:0] ethmac_writer_fifo_level = 2'd0;
reg ethmac_writer_fifo_replace = 1'd0;
reg ethmac_writer_fifo_produce = 1'd0;
reg ethmac_writer_fifo_consume = 1'd0;
reg ethmac_writer_fifo_wrport_adr = 1'd0;
wire [34:0] ethmac_writer_fifo_wrport_dat_r;
wire ethmac_writer_fifo_wrport_we;
wire [34:0] ethmac_writer_fifo_wrport_dat_w;
wire ethmac_writer_fifo_do_read;
wire ethmac_writer_fifo_rdport_adr;
wire [34:0] ethmac_writer_fifo_rdport_dat_r;
wire ethmac_writer_fifo_fifo_in_payload_slot;
wire [31:0] ethmac_writer_fifo_fifo_in_payload_length;
wire ethmac_writer_fifo_fifo_in_first;
wire ethmac_writer_fifo_fifo_in_last;
wire ethmac_writer_fifo_fifo_out_payload_slot;
wire [31:0] ethmac_writer_fifo_fifo_out_payload_length;
wire ethmac_writer_fifo_fifo_out_first;
wire ethmac_writer_fifo_fifo_out_last;
reg [8:0] ethmac_writer_memory0_adr = 9'd0;
wire [31:0] ethmac_writer_memory0_dat_r;
reg ethmac_writer_memory0_we = 1'd0;
reg [31:0] ethmac_writer_memory0_dat_w = 32'd0;
reg [8:0] ethmac_writer_memory1_adr = 9'd0;
wire [31:0] ethmac_writer_memory1_dat_r;
reg ethmac_writer_memory1_we = 1'd0;
reg [31:0] ethmac_writer_memory1_dat_w = 32'd0;
reg ethmac_reader_source_source_valid = 1'd0;
wire ethmac_reader_source_source_ready;
reg ethmac_reader_source_source_first = 1'd0;
reg ethmac_reader_source_source_last = 1'd0;
reg [31:0] ethmac_reader_source_source_payload_data = 32'd0;
reg [3:0] ethmac_reader_source_source_payload_last_be = 4'd0;
reg [3:0] ethmac_reader_source_source_payload_error = 4'd0;
wire ethmac_reader_start_re;
wire ethmac_reader_start_r;
reg ethmac_reader_start_w = 1'd0;
wire ethmac_reader_ready_status;
wire [1:0] ethmac_reader_level_status;
reg ethmac_reader_slot_storage_full = 1'd0;
wire ethmac_reader_slot_storage;
reg ethmac_reader_slot_re = 1'd0;
reg [10:0] ethmac_reader_length_storage_full = 11'd0;
wire [10:0] ethmac_reader_length_storage;
reg ethmac_reader_length_re = 1'd0;
wire ethmac_reader_irq;
wire ethmac_reader_done_status;
reg ethmac_reader_done_pending = 1'd0;
reg ethmac_reader_done_trigger = 1'd0;
reg ethmac_reader_done_clear = 1'd0;
wire ethmac_reader_eventmanager_status_re;
wire ethmac_reader_eventmanager_status_r;
wire ethmac_reader_eventmanager_status_w;
wire ethmac_reader_eventmanager_pending_re;
wire ethmac_reader_eventmanager_pending_r;
wire ethmac_reader_eventmanager_pending_w;
reg ethmac_reader_eventmanager_storage_full = 1'd0;
wire ethmac_reader_eventmanager_storage;
reg ethmac_reader_eventmanager_re = 1'd0;
wire ethmac_reader_fifo_sink_valid;
wire ethmac_reader_fifo_sink_ready;
reg ethmac_reader_fifo_sink_first = 1'd0;
reg ethmac_reader_fifo_sink_last = 1'd0;
wire ethmac_reader_fifo_sink_payload_slot;
wire [10:0] ethmac_reader_fifo_sink_payload_length;
wire ethmac_reader_fifo_source_valid;
reg ethmac_reader_fifo_source_ready = 1'd0;
wire ethmac_reader_fifo_source_first;
wire ethmac_reader_fifo_source_last;
wire ethmac_reader_fifo_source_payload_slot;
wire [10:0] ethmac_reader_fifo_source_payload_length;
wire ethmac_reader_fifo_syncfifo_we;
wire ethmac_reader_fifo_syncfifo_writable;
wire ethmac_reader_fifo_syncfifo_re;
wire ethmac_reader_fifo_syncfifo_readable;
wire [13:0] ethmac_reader_fifo_syncfifo_din;
wire [13:0] ethmac_reader_fifo_syncfifo_dout;
reg [1:0] ethmac_reader_fifo_level = 2'd0;
reg ethmac_reader_fifo_replace = 1'd0;
reg ethmac_reader_fifo_produce = 1'd0;
reg ethmac_reader_fifo_consume = 1'd0;
reg ethmac_reader_fifo_wrport_adr = 1'd0;
wire [13:0] ethmac_reader_fifo_wrport_dat_r;
wire ethmac_reader_fifo_wrport_we;
wire [13:0] ethmac_reader_fifo_wrport_dat_w;
wire ethmac_reader_fifo_do_read;
wire ethmac_reader_fifo_rdport_adr;
wire [13:0] ethmac_reader_fifo_rdport_dat_r;
wire ethmac_reader_fifo_fifo_in_payload_slot;
wire [10:0] ethmac_reader_fifo_fifo_in_payload_length;
wire ethmac_reader_fifo_fifo_in_first;
wire ethmac_reader_fifo_fifo_in_last;
wire ethmac_reader_fifo_fifo_out_payload_slot;
wire [10:0] ethmac_reader_fifo_fifo_out_payload_length;
wire ethmac_reader_fifo_fifo_out_first;
wire ethmac_reader_fifo_fifo_out_last;
reg [10:0] ethmac_reader_counter = 11'd0;
reg ethmac_reader_counter_reset = 1'd0;
reg ethmac_reader_counter_ce = 1'd0;
wire ethmac_reader_last;
reg ethmac_reader_last_d = 1'd0;
wire [8:0] ethmac_reader_memory0_adr;
wire [31:0] ethmac_reader_memory0_dat_r;
wire [8:0] ethmac_reader_memory1_adr;
wire [31:0] ethmac_reader_memory1_dat_r;
wire ethmac_ev_irq;
wire [29:0] ethmac_sram0_bus_adr0;
wire [31:0] ethmac_sram0_bus_dat_w0;
wire [31:0] ethmac_sram0_bus_dat_r0;
wire [3:0] ethmac_sram0_bus_sel0;
wire ethmac_sram0_bus_cyc0;
wire ethmac_sram0_bus_stb0;
reg ethmac_sram0_bus_ack0 = 1'd0;
wire ethmac_sram0_bus_we0;
wire [2:0] ethmac_sram0_bus_cti0;
wire [1:0] ethmac_sram0_bus_bte0;
reg ethmac_sram0_bus_err0 = 1'd0;
wire [8:0] ethmac_sram0_adr0;
wire [31:0] ethmac_sram0_dat_r0;
wire [29:0] ethmac_sram1_bus_adr0;
wire [31:0] ethmac_sram1_bus_dat_w0;
wire [31:0] ethmac_sram1_bus_dat_r0;
wire [3:0] ethmac_sram1_bus_sel0;
wire ethmac_sram1_bus_cyc0;
wire ethmac_sram1_bus_stb0;
reg ethmac_sram1_bus_ack0 = 1'd0;
wire ethmac_sram1_bus_we0;
wire [2:0] ethmac_sram1_bus_cti0;
wire [1:0] ethmac_sram1_bus_bte0;
reg ethmac_sram1_bus_err0 = 1'd0;
wire [8:0] ethmac_sram1_adr0;
wire [31:0] ethmac_sram1_dat_r0;
wire [29:0] ethmac_sram0_bus_adr1;
wire [31:0] ethmac_sram0_bus_dat_w1;
wire [31:0] ethmac_sram0_bus_dat_r1;
wire [3:0] ethmac_sram0_bus_sel1;
wire ethmac_sram0_bus_cyc1;
wire ethmac_sram0_bus_stb1;
reg ethmac_sram0_bus_ack1 = 1'd0;
wire ethmac_sram0_bus_we1;
wire [2:0] ethmac_sram0_bus_cti1;
wire [1:0] ethmac_sram0_bus_bte1;
reg ethmac_sram0_bus_err1 = 1'd0;
wire [8:0] ethmac_sram0_adr1;
wire [31:0] ethmac_sram0_dat_r1;
reg [3:0] ethmac_sram0_we = 4'd0;
wire [31:0] ethmac_sram0_dat_w;
wire [29:0] ethmac_sram1_bus_adr1;
wire [31:0] ethmac_sram1_bus_dat_w1;
wire [31:0] ethmac_sram1_bus_dat_r1;
wire [3:0] ethmac_sram1_bus_sel1;
wire ethmac_sram1_bus_cyc1;
wire ethmac_sram1_bus_stb1;
reg ethmac_sram1_bus_ack1 = 1'd0;
wire ethmac_sram1_bus_we1;
wire [2:0] ethmac_sram1_bus_cti1;
wire [1:0] ethmac_sram1_bus_bte1;
reg ethmac_sram1_bus_err1 = 1'd0;
wire [8:0] ethmac_sram1_adr1;
wire [31:0] ethmac_sram1_dat_r1;
reg [3:0] ethmac_sram1_we = 4'd0;
wire [31:0] ethmac_sram1_dat_w;
reg [3:0] ethmac_slave_sel = 4'd0;
reg [3:0] ethmac_slave_sel_r = 4'd0;
wire litedramcrossbar_cmd_valid;
wire litedramcrossbar_cmd_ready;
wire litedramcrossbar_cmd_payload_we;
wire [24:0] litedramcrossbar_cmd_payload_adr;
wire litedramcrossbar_wdata_valid;
wire litedramcrossbar_wdata_ready;
wire [127:0] litedramcrossbar_wdata_payload_data;
wire [15:0] litedramcrossbar_wdata_payload_we;
wire litedramcrossbar_rdata_valid;
wire [127:0] litedramcrossbar_rdata_payload_data;
wire edid_status;
reg edid_storage_full = 1'd0;
wire edid_storage;
reg edid_re = 1'd0;
wire edid_scl_raw;
reg edid_sda_i = 1'd0;
wire edid_sda_raw;
reg edid_sda_drv = 1'd0;
reg edid_sda_drv_reg = 1'd0;
wire edid_sda_i_async;
wire edid_sda_o;
reg edid_scl_i = 1'd0;
reg [5:0] edid_samp_count = 6'd0;
reg edid_samp_carry = 1'd0;
reg edid_scl_r = 1'd0;
reg edid_sda_r = 1'd0;
wire edid_scl_rising;
wire edid_sda_rising;
wire edid_sda_falling;
wire edid_start;
reg [7:0] edid_din = 8'd0;
reg [3:0] edid_counter = 4'd0;
reg edid_is_read = 1'd0;
reg edid_update_is_read = 1'd0;
reg [6:0] edid_offset_counter = 7'd0;
reg edid_oc_load = 1'd0;
reg edid_oc_inc = 1'd0;
wire [6:0] edid_adr;
wire [7:0] edid_dat_r;
reg edid_data_bit = 1'd0;
reg edid_zero_drv = 1'd0;
reg edid_data_drv = 1'd0;
reg edid_data_drv_en = 1'd0;
reg edid_data_drv_stop = 1'd0;
reg mmcm_reset_storage_full = 1'd1;
wire mmcm_reset_storage;
reg mmcm_reset_re = 1'd0;
wire locked_status;
wire mmcm_read_re;
wire mmcm_read_r;
reg mmcm_read_w = 1'd0;
wire mmcm_write_re;
wire mmcm_write_r;
reg mmcm_write_w = 1'd0;
reg mmcm_drdy_status = 1'd0;
reg [6:0] mmcm_adr_storage_full = 7'd0;
wire [6:0] mmcm_adr_storage;
reg mmcm_adr_re = 1'd0;
reg [15:0] mmcm_dat_w_storage_full = 16'd0;
wire [15:0] mmcm_dat_w_storage;
reg mmcm_dat_w_re = 1'd0;
wire [15:0] mmcm_dat_r_status;
wire locked;
wire hdmi_in0_pix_clk;
wire hdmi_in0_pix_rst;
wire pix1p25x_clk;
wire pix1p25x_rst;
wire hdmi_in0_pix5x_clk;
wire clk_input;
wire clk_input_bufg;
wire mmcm_fb;
wire mmcm_locked;
wire mmcm_clk0;
wire mmcm_clk1;
wire mmcm_clk2;
wire mmcm_drdy;
wire [9:0] s7datacapture0_d;
wire s7datacapture0_dly_ctl_re;
wire [4:0] s7datacapture0_dly_ctl_r;
reg [4:0] s7datacapture0_dly_ctl_w = 5'd0;
wire [1:0] s7datacapture0_status;
wire s7datacapture0_phase_reset_re;
wire s7datacapture0_phase_reset_r;
reg s7datacapture0_phase_reset_w = 1'd0;
wire s7datacapture0_serdes_m_i_nodelay;
wire s7datacapture0_serdes_s_i_nodelay;
wire s7datacapture0_delay_rst;
wire s7datacapture0_delay_master_inc;
wire s7datacapture0_delay_master_ce;
wire s7datacapture0_delay_slave_inc;
wire s7datacapture0_delay_slave_ce;
wire s7datacapture0_serdes_m_i_delayed;
wire [7:0] s7datacapture0_serdes_m_q;
wire [7:0] s7datacapture0_serdes_m_d;
wire s7datacapture0_serdes_s_i_delayed;
wire [7:0] s7datacapture0_serdes_s_q;
wire [7:0] s7datacapture0_serdes_s_d;
wire [7:0] s7datacapture0_gearbox_i;
reg [9:0] s7datacapture0_gearbox_o = 10'd0;
wire s7datacapture0_gearbox_rst;
wire data0_cap_write_clk;
wire data0_cap_write_rst;
wire data0_cap_read_clk;
wire data0_cap_read_rst;
reg [79:0] s7datacapture0_gearbox_storage = 80'd0;
reg [3:0] s7datacapture0_gearbox_wrpointer = 4'd5;
reg [2:0] s7datacapture0_gearbox_rdpointer = 3'd0;
wire [7:0] s7datacapture0_mdata;
wire [7:0] s7datacapture0_sdata;
wire s7datacapture0_inc;
wire s7datacapture0_dec;
wire s7datacapture0_transition;
reg [7:0] s7datacapture0_mdata_d = 8'd0;
reg [7:0] s7datacapture0_lateness = 8'd128;
wire s7datacapture0_too_late;
wire s7datacapture0_too_early;
wire s7datacapture0_reset_lateness;
wire s7datacapture0_do_delay_rst_i;
wire s7datacapture0_do_delay_rst_o;
reg s7datacapture0_do_delay_rst_toggle_i = 1'd0;
wire s7datacapture0_do_delay_rst_toggle_o;
reg s7datacapture0_do_delay_rst_toggle_o_r = 1'd0;
wire s7datacapture0_do_delay_master_inc_i;
wire s7datacapture0_do_delay_master_inc_o;
reg s7datacapture0_do_delay_master_inc_toggle_i = 1'd0;
wire s7datacapture0_do_delay_master_inc_toggle_o;
reg s7datacapture0_do_delay_master_inc_toggle_o_r = 1'd0;
wire s7datacapture0_do_delay_master_dec_i;
wire s7datacapture0_do_delay_master_dec_o;
reg s7datacapture0_do_delay_master_dec_toggle_i = 1'd0;
wire s7datacapture0_do_delay_master_dec_toggle_o;
reg s7datacapture0_do_delay_master_dec_toggle_o_r = 1'd0;
wire s7datacapture0_do_delay_slave_inc_i;
wire s7datacapture0_do_delay_slave_inc_o;
reg s7datacapture0_do_delay_slave_inc_toggle_i = 1'd0;
wire s7datacapture0_do_delay_slave_inc_toggle_o;
reg s7datacapture0_do_delay_slave_inc_toggle_o_r = 1'd0;
wire s7datacapture0_do_delay_slave_dec_i;
wire s7datacapture0_do_delay_slave_dec_o;
reg s7datacapture0_do_delay_slave_dec_toggle_i = 1'd0;
wire s7datacapture0_do_delay_slave_dec_toggle_o;
reg s7datacapture0_do_delay_slave_dec_toggle_o_r = 1'd0;
wire s7datacapture0_do_reset_lateness_i;
wire s7datacapture0_do_reset_lateness_o;
reg s7datacapture0_do_reset_lateness_toggle_i = 1'd0;
wire s7datacapture0_do_reset_lateness_toggle_o;
reg s7datacapture0_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] charsync0_raw_data;
reg charsync0_synced = 1'd0;
reg [9:0] charsync0_data = 10'd0;
wire charsync0_char_synced_status;
wire [3:0] charsync0_ctl_pos_status;
reg [9:0] charsync0_raw_data1 = 10'd0;
wire [19:0] charsync0_raw;
reg charsync0_found_control = 1'd0;
reg [3:0] charsync0_control_position = 4'd0;
reg [2:0] charsync0_control_counter = 3'd0;
reg [3:0] charsync0_previous_control_position = 4'd0;
reg [3:0] charsync0_word_sel = 4'd0;
wire [9:0] wer0_data;
wire wer0_update_re;
wire wer0_update_r;
reg wer0_update_w = 1'd0;
reg [23:0] wer0_status = 24'd0;
reg [8:0] wer0_data_r = 9'd0;
reg [7:0] wer0_transitions = 8'd0;
reg [3:0] wer0_transition_count = 4'd0;
reg wer0_is_control = 1'd0;
reg wer0_is_error = 1'd0;
reg [23:0] wer0_period_counter = 24'd0;
reg wer0_period_done = 1'd0;
reg [23:0] wer0_wer_counter = 24'd0;
reg [23:0] wer0_wer_counter_r = 24'd0;
reg wer0_wer_counter_r_updated = 1'd0;
reg [23:0] wer0_wer_counter_sys = 24'd0;
wire wer0_i;
wire wer0_o;
reg wer0_toggle_i = 1'd0;
wire wer0_toggle_o;
reg wer0_toggle_o_r = 1'd0;
wire decoding0_valid_i;
wire [9:0] decoding0_input;
reg decoding0_valid_o = 1'd0;
reg [7:0] decoding0_output_d = 8'd0;
reg [1:0] decoding0_output_c = 2'd0;
reg decoding0_output_de = 1'd0;
wire [9:0] s7datacapture1_d;
wire s7datacapture1_dly_ctl_re;
wire [4:0] s7datacapture1_dly_ctl_r;
reg [4:0] s7datacapture1_dly_ctl_w = 5'd0;
wire [1:0] s7datacapture1_status;
wire s7datacapture1_phase_reset_re;
wire s7datacapture1_phase_reset_r;
reg s7datacapture1_phase_reset_w = 1'd0;
wire s7datacapture1_serdes_m_i_nodelay;
wire s7datacapture1_serdes_s_i_nodelay;
wire s7datacapture1_delay_rst;
wire s7datacapture1_delay_master_inc;
wire s7datacapture1_delay_master_ce;
wire s7datacapture1_delay_slave_inc;
wire s7datacapture1_delay_slave_ce;
wire s7datacapture1_serdes_m_i_delayed;
wire [7:0] s7datacapture1_serdes_m_q;
wire [7:0] s7datacapture1_serdes_m_d;
wire s7datacapture1_serdes_s_i_delayed;
wire [7:0] s7datacapture1_serdes_s_q;
wire [7:0] s7datacapture1_serdes_s_d;
wire [7:0] s7datacapture1_gearbox_i;
reg [9:0] s7datacapture1_gearbox_o = 10'd0;
wire s7datacapture1_gearbox_rst;
wire data1_cap_write_clk;
wire data1_cap_write_rst;
wire data1_cap_read_clk;
wire data1_cap_read_rst;
reg [79:0] s7datacapture1_gearbox_storage = 80'd0;
reg [3:0] s7datacapture1_gearbox_wrpointer = 4'd5;
reg [2:0] s7datacapture1_gearbox_rdpointer = 3'd0;
wire [7:0] s7datacapture1_mdata;
wire [7:0] s7datacapture1_sdata;
wire s7datacapture1_inc;
wire s7datacapture1_dec;
wire s7datacapture1_transition;
reg [7:0] s7datacapture1_mdata_d = 8'd0;
reg [7:0] s7datacapture1_lateness = 8'd128;
wire s7datacapture1_too_late;
wire s7datacapture1_too_early;
wire s7datacapture1_reset_lateness;
wire s7datacapture1_do_delay_rst_i;
wire s7datacapture1_do_delay_rst_o;
reg s7datacapture1_do_delay_rst_toggle_i = 1'd0;
wire s7datacapture1_do_delay_rst_toggle_o;
reg s7datacapture1_do_delay_rst_toggle_o_r = 1'd0;
wire s7datacapture1_do_delay_master_inc_i;
wire s7datacapture1_do_delay_master_inc_o;
reg s7datacapture1_do_delay_master_inc_toggle_i = 1'd0;
wire s7datacapture1_do_delay_master_inc_toggle_o;
reg s7datacapture1_do_delay_master_inc_toggle_o_r = 1'd0;
wire s7datacapture1_do_delay_master_dec_i;
wire s7datacapture1_do_delay_master_dec_o;
reg s7datacapture1_do_delay_master_dec_toggle_i = 1'd0;
wire s7datacapture1_do_delay_master_dec_toggle_o;
reg s7datacapture1_do_delay_master_dec_toggle_o_r = 1'd0;
wire s7datacapture1_do_delay_slave_inc_i;
wire s7datacapture1_do_delay_slave_inc_o;
reg s7datacapture1_do_delay_slave_inc_toggle_i = 1'd0;
wire s7datacapture1_do_delay_slave_inc_toggle_o;
reg s7datacapture1_do_delay_slave_inc_toggle_o_r = 1'd0;
wire s7datacapture1_do_delay_slave_dec_i;
wire s7datacapture1_do_delay_slave_dec_o;
reg s7datacapture1_do_delay_slave_dec_toggle_i = 1'd0;
wire s7datacapture1_do_delay_slave_dec_toggle_o;
reg s7datacapture1_do_delay_slave_dec_toggle_o_r = 1'd0;
wire s7datacapture1_do_reset_lateness_i;
wire s7datacapture1_do_reset_lateness_o;
reg s7datacapture1_do_reset_lateness_toggle_i = 1'd0;
wire s7datacapture1_do_reset_lateness_toggle_o;
reg s7datacapture1_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] charsync1_raw_data;
reg charsync1_synced = 1'd0;
reg [9:0] charsync1_data = 10'd0;
wire charsync1_char_synced_status;
wire [3:0] charsync1_ctl_pos_status;
reg [9:0] charsync1_raw_data1 = 10'd0;
wire [19:0] charsync1_raw;
reg charsync1_found_control = 1'd0;
reg [3:0] charsync1_control_position = 4'd0;
reg [2:0] charsync1_control_counter = 3'd0;
reg [3:0] charsync1_previous_control_position = 4'd0;
reg [3:0] charsync1_word_sel = 4'd0;
wire [9:0] wer1_data;
wire wer1_update_re;
wire wer1_update_r;
reg wer1_update_w = 1'd0;
reg [23:0] wer1_status = 24'd0;
reg [8:0] wer1_data_r = 9'd0;
reg [7:0] wer1_transitions = 8'd0;
reg [3:0] wer1_transition_count = 4'd0;
reg wer1_is_control = 1'd0;
reg wer1_is_error = 1'd0;
reg [23:0] wer1_period_counter = 24'd0;
reg wer1_period_done = 1'd0;
reg [23:0] wer1_wer_counter = 24'd0;
reg [23:0] wer1_wer_counter_r = 24'd0;
reg wer1_wer_counter_r_updated = 1'd0;
reg [23:0] wer1_wer_counter_sys = 24'd0;
wire wer1_i;
wire wer1_o;
reg wer1_toggle_i = 1'd0;
wire wer1_toggle_o;
reg wer1_toggle_o_r = 1'd0;
wire decoding1_valid_i;
wire [9:0] decoding1_input;
reg decoding1_valid_o = 1'd0;
reg [7:0] decoding1_output_d = 8'd0;
reg [1:0] decoding1_output_c = 2'd0;
reg decoding1_output_de = 1'd0;
wire [9:0] s7datacapture2_d;
wire s7datacapture2_dly_ctl_re;
wire [4:0] s7datacapture2_dly_ctl_r;
reg [4:0] s7datacapture2_dly_ctl_w = 5'd0;
wire [1:0] s7datacapture2_status;
wire s7datacapture2_phase_reset_re;
wire s7datacapture2_phase_reset_r;
reg s7datacapture2_phase_reset_w = 1'd0;
wire s7datacapture2_serdes_m_i_nodelay;
wire s7datacapture2_serdes_s_i_nodelay;
wire s7datacapture2_delay_rst;
wire s7datacapture2_delay_master_inc;
wire s7datacapture2_delay_master_ce;
wire s7datacapture2_delay_slave_inc;
wire s7datacapture2_delay_slave_ce;
wire s7datacapture2_serdes_m_i_delayed;
wire [7:0] s7datacapture2_serdes_m_q;
wire [7:0] s7datacapture2_serdes_m_d;
wire s7datacapture2_serdes_s_i_delayed;
wire [7:0] s7datacapture2_serdes_s_q;
wire [7:0] s7datacapture2_serdes_s_d;
wire [7:0] s7datacapture2_gearbox_i;
reg [9:0] s7datacapture2_gearbox_o = 10'd0;
wire s7datacapture2_gearbox_rst;
wire data2_cap_write_clk;
wire data2_cap_write_rst;
wire data2_cap_read_clk;
wire data2_cap_read_rst;
reg [79:0] s7datacapture2_gearbox_storage = 80'd0;
reg [3:0] s7datacapture2_gearbox_wrpointer = 4'd5;
reg [2:0] s7datacapture2_gearbox_rdpointer = 3'd0;
wire [7:0] s7datacapture2_mdata;
wire [7:0] s7datacapture2_sdata;
wire s7datacapture2_inc;
wire s7datacapture2_dec;
wire s7datacapture2_transition;
reg [7:0] s7datacapture2_mdata_d = 8'd0;
reg [7:0] s7datacapture2_lateness = 8'd128;
wire s7datacapture2_too_late;
wire s7datacapture2_too_early;
wire s7datacapture2_reset_lateness;
wire s7datacapture2_do_delay_rst_i;
wire s7datacapture2_do_delay_rst_o;
reg s7datacapture2_do_delay_rst_toggle_i = 1'd0;
wire s7datacapture2_do_delay_rst_toggle_o;
reg s7datacapture2_do_delay_rst_toggle_o_r = 1'd0;
wire s7datacapture2_do_delay_master_inc_i;
wire s7datacapture2_do_delay_master_inc_o;
reg s7datacapture2_do_delay_master_inc_toggle_i = 1'd0;
wire s7datacapture2_do_delay_master_inc_toggle_o;
reg s7datacapture2_do_delay_master_inc_toggle_o_r = 1'd0;
wire s7datacapture2_do_delay_master_dec_i;
wire s7datacapture2_do_delay_master_dec_o;
reg s7datacapture2_do_delay_master_dec_toggle_i = 1'd0;
wire s7datacapture2_do_delay_master_dec_toggle_o;
reg s7datacapture2_do_delay_master_dec_toggle_o_r = 1'd0;
wire s7datacapture2_do_delay_slave_inc_i;
wire s7datacapture2_do_delay_slave_inc_o;
reg s7datacapture2_do_delay_slave_inc_toggle_i = 1'd0;
wire s7datacapture2_do_delay_slave_inc_toggle_o;
reg s7datacapture2_do_delay_slave_inc_toggle_o_r = 1'd0;
wire s7datacapture2_do_delay_slave_dec_i;
wire s7datacapture2_do_delay_slave_dec_o;
reg s7datacapture2_do_delay_slave_dec_toggle_i = 1'd0;
wire s7datacapture2_do_delay_slave_dec_toggle_o;
reg s7datacapture2_do_delay_slave_dec_toggle_o_r = 1'd0;
wire s7datacapture2_do_reset_lateness_i;
wire s7datacapture2_do_reset_lateness_o;
reg s7datacapture2_do_reset_lateness_toggle_i = 1'd0;
wire s7datacapture2_do_reset_lateness_toggle_o;
reg s7datacapture2_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] charsync2_raw_data;
reg charsync2_synced = 1'd0;
reg [9:0] charsync2_data = 10'd0;
wire charsync2_char_synced_status;
wire [3:0] charsync2_ctl_pos_status;
reg [9:0] charsync2_raw_data1 = 10'd0;
wire [19:0] charsync2_raw;
reg charsync2_found_control = 1'd0;
reg [3:0] charsync2_control_position = 4'd0;
reg [2:0] charsync2_control_counter = 3'd0;
reg [3:0] charsync2_previous_control_position = 4'd0;
reg [3:0] charsync2_word_sel = 4'd0;
wire [9:0] wer2_data;
wire wer2_update_re;
wire wer2_update_r;
reg wer2_update_w = 1'd0;
reg [23:0] wer2_status = 24'd0;
reg [8:0] wer2_data_r = 9'd0;
reg [7:0] wer2_transitions = 8'd0;
reg [3:0] wer2_transition_count = 4'd0;
reg wer2_is_control = 1'd0;
reg wer2_is_error = 1'd0;
reg [23:0] wer2_period_counter = 24'd0;
reg wer2_period_done = 1'd0;
reg [23:0] wer2_wer_counter = 24'd0;
reg [23:0] wer2_wer_counter_r = 24'd0;
reg wer2_wer_counter_r_updated = 1'd0;
reg [23:0] wer2_wer_counter_sys = 24'd0;
wire wer2_i;
wire wer2_o;
reg wer2_toggle_i = 1'd0;
wire wer2_toggle_o;
reg wer2_toggle_o_r = 1'd0;
wire decoding2_valid_i;
wire [9:0] decoding2_input;
reg decoding2_valid_o = 1'd0;
reg [7:0] decoding2_output_d = 8'd0;
reg [1:0] decoding2_output_c = 2'd0;
reg decoding2_output_de = 1'd0;
wire chansync_valid_i;
reg chansync_chan_synced = 1'd0;
wire chansync_status;
wire chansync_all_control;
wire [7:0] chansync_data_in0_d;
wire [1:0] chansync_data_in0_c;
wire chansync_data_in0_de;
wire [7:0] chansync_data_out0_d;
wire [1:0] chansync_data_out0_c;
wire chansync_data_out0_de;
wire [10:0] chansync_syncbuffer0_din;
wire [10:0] chansync_syncbuffer0_dout;
wire chansync_syncbuffer0_re;
reg [2:0] chansync_syncbuffer0_produce = 3'd0;
reg [2:0] chansync_syncbuffer0_consume = 3'd0;
wire [2:0] chansync_syncbuffer0_wrport_adr;
wire [10:0] chansync_syncbuffer0_wrport_dat_r;
wire chansync_syncbuffer0_wrport_we;
wire [10:0] chansync_syncbuffer0_wrport_dat_w;
wire [2:0] chansync_syncbuffer0_rdport_adr;
wire [10:0] chansync_syncbuffer0_rdport_dat_r;
wire chansync_is_control0;
wire [7:0] chansync_data_in1_d;
wire [1:0] chansync_data_in1_c;
wire chansync_data_in1_de;
wire [7:0] chansync_data_out1_d;
wire [1:0] chansync_data_out1_c;
wire chansync_data_out1_de;
wire [10:0] chansync_syncbuffer1_din;
wire [10:0] chansync_syncbuffer1_dout;
wire chansync_syncbuffer1_re;
reg [2:0] chansync_syncbuffer1_produce = 3'd0;
reg [2:0] chansync_syncbuffer1_consume = 3'd0;
wire [2:0] chansync_syncbuffer1_wrport_adr;
wire [10:0] chansync_syncbuffer1_wrport_dat_r;
wire chansync_syncbuffer1_wrport_we;
wire [10:0] chansync_syncbuffer1_wrport_dat_w;
wire [2:0] chansync_syncbuffer1_rdport_adr;
wire [10:0] chansync_syncbuffer1_rdport_dat_r;
wire chansync_is_control1;
wire [7:0] chansync_data_in2_d;
wire [1:0] chansync_data_in2_c;
wire chansync_data_in2_de;
wire [7:0] chansync_data_out2_d;
wire [1:0] chansync_data_out2_c;
wire chansync_data_out2_de;
wire [10:0] chansync_syncbuffer2_din;
wire [10:0] chansync_syncbuffer2_dout;
wire chansync_syncbuffer2_re;
reg [2:0] chansync_syncbuffer2_produce = 3'd0;
reg [2:0] chansync_syncbuffer2_consume = 3'd0;
wire [2:0] chansync_syncbuffer2_wrport_adr;
wire [10:0] chansync_syncbuffer2_wrport_dat_r;
wire chansync_syncbuffer2_wrport_we;
wire [10:0] chansync_syncbuffer2_wrport_dat_w;
wire [2:0] chansync_syncbuffer2_rdport_adr;
wire [10:0] chansync_syncbuffer2_rdport_dat_r;
wire chansync_is_control2;
wire chansync_some_control;
wire syncpol_valid_i;
wire [7:0] syncpol_data_in0_d;
wire [1:0] syncpol_data_in0_c;
wire syncpol_data_in0_de;
wire [7:0] syncpol_data_in1_d;
wire [1:0] syncpol_data_in1_c;
wire syncpol_data_in1_de;
wire [7:0] syncpol_data_in2_d;
wire [1:0] syncpol_data_in2_c;
wire syncpol_data_in2_de;
reg syncpol_valid_o = 1'd0;
wire syncpol_de;
wire syncpol_hsync;
wire syncpol_vsync;
reg [7:0] syncpol_r = 8'd0;
reg [7:0] syncpol_g = 8'd0;
reg [7:0] syncpol_b = 8'd0;
reg syncpol_de_r = 1'd0;
reg [1:0] syncpol_c_polarity = 2'd0;
reg [1:0] syncpol_c_out = 2'd0;
wire resdetection_valid_i;
wire resdetection_vsync;
wire resdetection_de;
wire [10:0] resdetection_hres_status;
wire [10:0] resdetection_vres_status;
reg resdetection_de_r = 1'd0;
wire resdetection_pn_de;
reg [10:0] resdetection_hcounter = 11'd0;
reg [10:0] resdetection_hcounter_st = 11'd0;
reg resdetection_vsync_r = 1'd0;
wire resdetection_p_vsync;
reg [10:0] resdetection_vcounter = 11'd0;
reg [10:0] resdetection_vcounter_st = 11'd0;
wire frame_valid_i;
wire frame_vsync;
wire frame_de;
wire [7:0] frame_r;
wire [7:0] frame_g;
wire [7:0] frame_b;
wire frame_frame_valid;
wire frame_frame_ready;
wire frame_frame_first;
wire frame_frame_last;
wire frame_frame_payload_sof;
wire [127:0] frame_frame_payload_pixels;
wire frame_busy;
wire frame_overflow_re;
wire frame_overflow_r;
wire frame_overflow_w;
reg frame_de_r = 1'd0;
wire frame_rgb2ycbcr_sink_valid;
wire frame_rgb2ycbcr_sink_ready;
reg frame_rgb2ycbcr_sink_first = 1'd0;
reg frame_rgb2ycbcr_sink_last = 1'd0;
wire [7:0] frame_rgb2ycbcr_sink_payload_r;
wire [7:0] frame_rgb2ycbcr_sink_payload_g;
wire [7:0] frame_rgb2ycbcr_sink_payload_b;
wire frame_rgb2ycbcr_source_valid;
wire frame_rgb2ycbcr_source_ready;
wire frame_rgb2ycbcr_source_first;
wire frame_rgb2ycbcr_source_last;
wire [7:0] frame_rgb2ycbcr_source_payload_y;
wire [7:0] frame_rgb2ycbcr_source_payload_cb;
wire [7:0] frame_rgb2ycbcr_source_payload_cr;
wire [7:0] frame_rgb2ycbcr_sink_r;
wire [7:0] frame_rgb2ycbcr_sink_g;
wire [7:0] frame_rgb2ycbcr_sink_b;
reg [7:0] frame_rgb2ycbcr_source_y = 8'd0;
reg [7:0] frame_rgb2ycbcr_source_cb = 8'd0;
reg [7:0] frame_rgb2ycbcr_source_cr = 8'd0;
reg [7:0] frame_rgb2ycbcr_record0_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record0_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record0_rgb_n_b = 8'd0;
reg [7:0] frame_rgb2ycbcr_record1_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record1_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record1_rgb_n_b = 8'd0;
reg [7:0] frame_rgb2ycbcr_record2_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record2_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record2_rgb_n_b = 8'd0;
reg [7:0] frame_rgb2ycbcr_record3_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record3_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record3_rgb_n_b = 8'd0;
reg [7:0] frame_rgb2ycbcr_record4_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record4_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record4_rgb_n_b = 8'd0;
reg [7:0] frame_rgb2ycbcr_record5_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record5_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record5_rgb_n_b = 8'd0;
reg [7:0] frame_rgb2ycbcr_record6_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record6_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record6_rgb_n_b = 8'd0;
reg [7:0] frame_rgb2ycbcr_record7_rgb_n_r = 8'd0;
reg [7:0] frame_rgb2ycbcr_record7_rgb_n_g = 8'd0;
reg [7:0] frame_rgb2ycbcr_record7_rgb_n_b = 8'd0;
reg signed [8:0] frame_rgb2ycbcr_r_minus_g = 9'sd512;
reg signed [8:0] frame_rgb2ycbcr_b_minus_g = 9'sd512;
reg signed [16:0] frame_rgb2ycbcr_ca_mult_rg = 17'sd131072;
reg signed [16:0] frame_rgb2ycbcr_cb_mult_bg = 17'sd131072;
reg signed [24:0] frame_rgb2ycbcr_carg_plus_cbbg = 25'sd33554432;
reg signed [10:0] frame_rgb2ycbcr_yraw = 11'sd2048;
reg signed [11:0] frame_rgb2ycbcr_b_minus_yraw = 12'sd4096;
reg signed [11:0] frame_rgb2ycbcr_r_minus_yraw = 12'sd4096;
reg signed [10:0] frame_rgb2ycbcr_yraw_r0 = 11'sd2048;
reg signed [19:0] frame_rgb2ycbcr_cc_mult_ryraw = 20'sd1048576;
reg signed [19:0] frame_rgb2ycbcr_cd_mult_byraw = 20'sd1048576;
reg signed [10:0] frame_rgb2ycbcr_yraw_r1 = 11'sd2048;
reg signed [10:0] frame_rgb2ycbcr_y = 11'sd2048;
reg signed [11:0] frame_rgb2ycbcr_cb = 12'sd4096;
reg signed [11:0] frame_rgb2ycbcr_cr = 12'sd4096;
wire frame_rgb2ycbcr_ce;
wire frame_rgb2ycbcr_pipe_ce;
wire frame_rgb2ycbcr_busy;
reg frame_rgb2ycbcr_valid_n0 = 1'd0;
reg frame_rgb2ycbcr_valid_n1 = 1'd0;
reg frame_rgb2ycbcr_valid_n2 = 1'd0;
reg frame_rgb2ycbcr_valid_n3 = 1'd0;
reg frame_rgb2ycbcr_valid_n4 = 1'd0;
reg frame_rgb2ycbcr_valid_n5 = 1'd0;
reg frame_rgb2ycbcr_valid_n6 = 1'd0;
reg frame_rgb2ycbcr_valid_n7 = 1'd0;
reg frame_rgb2ycbcr_first_n0 = 1'd0;
reg frame_rgb2ycbcr_last_n0 = 1'd0;
reg frame_rgb2ycbcr_first_n1 = 1'd0;
reg frame_rgb2ycbcr_last_n1 = 1'd0;
reg frame_rgb2ycbcr_first_n2 = 1'd0;
reg frame_rgb2ycbcr_last_n2 = 1'd0;
reg frame_rgb2ycbcr_first_n3 = 1'd0;
reg frame_rgb2ycbcr_last_n3 = 1'd0;
reg frame_rgb2ycbcr_first_n4 = 1'd0;
reg frame_rgb2ycbcr_last_n4 = 1'd0;
reg frame_rgb2ycbcr_first_n5 = 1'd0;
reg frame_rgb2ycbcr_last_n5 = 1'd0;
reg frame_rgb2ycbcr_first_n6 = 1'd0;
reg frame_rgb2ycbcr_last_n6 = 1'd0;
reg frame_rgb2ycbcr_first_n7 = 1'd0;
reg frame_rgb2ycbcr_last_n7 = 1'd0;
wire frame_chroma_downsampler_sink_valid;
wire frame_chroma_downsampler_sink_ready;
wire frame_chroma_downsampler_sink_first;
wire frame_chroma_downsampler_sink_last;
wire [7:0] frame_chroma_downsampler_sink_payload_y;
wire [7:0] frame_chroma_downsampler_sink_payload_cb;
wire [7:0] frame_chroma_downsampler_sink_payload_cr;
wire frame_chroma_downsampler_source_valid;
wire frame_chroma_downsampler_source_ready;
wire frame_chroma_downsampler_source_first;
wire frame_chroma_downsampler_source_last;
wire [7:0] frame_chroma_downsampler_source_payload_y;
wire [7:0] frame_chroma_downsampler_source_payload_cb_cr;
wire [7:0] frame_chroma_downsampler_sink_y;
wire [7:0] frame_chroma_downsampler_sink_cb;
wire [7:0] frame_chroma_downsampler_sink_cr;
reg [7:0] frame_chroma_downsampler_source_y = 8'd0;
reg [7:0] frame_chroma_downsampler_source_cb_cr = 8'd0;
wire frame_chroma_downsampler_first;
reg [7:0] frame_chroma_downsampler_record0_ycbcr_n_y = 8'd0;
reg [7:0] frame_chroma_downsampler_record0_ycbcr_n_cb = 8'd0;
reg [7:0] frame_chroma_downsampler_record0_ycbcr_n_cr = 8'd0;
reg [7:0] frame_chroma_downsampler_record1_ycbcr_n_y = 8'd0;
reg [7:0] frame_chroma_downsampler_record1_ycbcr_n_cb = 8'd0;
reg [7:0] frame_chroma_downsampler_record1_ycbcr_n_cr = 8'd0;
reg [7:0] frame_chroma_downsampler_record2_ycbcr_n_y = 8'd0;
reg [7:0] frame_chroma_downsampler_record2_ycbcr_n_cb = 8'd0;
reg [7:0] frame_chroma_downsampler_record2_ycbcr_n_cr = 8'd0;
reg frame_chroma_downsampler_parity = 1'd0;
reg [8:0] frame_chroma_downsampler_cb_sum = 9'd0;
reg [8:0] frame_chroma_downsampler_cr_sum = 9'd0;
wire [7:0] frame_chroma_downsampler_cb_mean;
wire [7:0] frame_chroma_downsampler_cr_mean;
wire frame_chroma_downsampler_ce;
wire frame_chroma_downsampler_pipe_ce;
wire frame_chroma_downsampler_busy;
reg frame_chroma_downsampler_valid_n0 = 1'd0;
reg frame_chroma_downsampler_valid_n1 = 1'd0;
reg frame_chroma_downsampler_valid_n2 = 1'd0;
reg frame_chroma_downsampler_first_n0 = 1'd0;
reg frame_chroma_downsampler_last_n0 = 1'd0;
reg frame_chroma_downsampler_first_n1 = 1'd0;
reg frame_chroma_downsampler_last_n1 = 1'd0;
reg frame_chroma_downsampler_first_n2 = 1'd0;
reg frame_chroma_downsampler_last_n2 = 1'd0;
reg frame_next_de0 = 1'd0;
reg frame_next_vsync0 = 1'd0;
reg frame_next_de1 = 1'd0;
reg frame_next_vsync1 = 1'd0;
reg frame_next_de2 = 1'd0;
reg frame_next_vsync2 = 1'd0;
reg frame_next_de3 = 1'd0;
reg frame_next_vsync3 = 1'd0;
reg frame_next_de4 = 1'd0;
reg frame_next_vsync4 = 1'd0;
reg frame_next_de5 = 1'd0;
reg frame_next_vsync5 = 1'd0;
reg frame_next_de6 = 1'd0;
reg frame_next_vsync6 = 1'd0;
reg frame_next_de7 = 1'd0;
reg frame_next_vsync7 = 1'd0;
reg frame_next_de8 = 1'd0;
reg frame_next_vsync8 = 1'd0;
reg frame_next_de9 = 1'd0;
reg frame_next_vsync9 = 1'd0;
reg frame_next_de10 = 1'd0;
reg frame_next_vsync10 = 1'd0;
reg frame_vsync_r = 1'd0;
wire frame_new_frame;
reg [127:0] frame_cur_word = 128'd0;
reg frame_cur_word_valid = 1'd0;
wire [15:0] frame_encoded_pixel;
reg [2:0] frame_pack_counter = 3'd0;
wire frame_fifo_sink_valid;
wire frame_fifo_sink_ready;
reg frame_fifo_sink_first = 1'd0;
reg frame_fifo_sink_last = 1'd0;
reg frame_fifo_sink_payload_sof = 1'd0;
wire [127:0] frame_fifo_sink_payload_pixels;
wire frame_fifo_source_valid;
wire frame_fifo_source_ready;
wire frame_fifo_source_first;
wire frame_fifo_source_last;
wire frame_fifo_source_payload_sof;
wire [127:0] frame_fifo_source_payload_pixels;
wire frame_fifo_asyncfifo_we;
wire frame_fifo_asyncfifo_writable;
wire frame_fifo_asyncfifo_re;
wire frame_fifo_asyncfifo_readable;
wire [130:0] frame_fifo_asyncfifo_din;
wire [130:0] frame_fifo_asyncfifo_dout;
wire frame_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [9:0] frame_fifo_graycounter0_q = 10'd0;
wire [9:0] frame_fifo_graycounter0_q_next;
reg [9:0] frame_fifo_graycounter0_q_binary = 10'd0;
reg [9:0] frame_fifo_graycounter0_q_next_binary = 10'd0;
wire frame_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [9:0] frame_fifo_graycounter1_q = 10'd0;
wire [9:0] frame_fifo_graycounter1_q_next;
reg [9:0] frame_fifo_graycounter1_q_binary = 10'd0;
reg [9:0] frame_fifo_graycounter1_q_next_binary = 10'd0;
wire [9:0] frame_fifo_produce_rdomain;
wire [9:0] frame_fifo_consume_wdomain;
wire [8:0] frame_fifo_wrport_adr;
wire [130:0] frame_fifo_wrport_dat_r;
wire frame_fifo_wrport_we;
wire [130:0] frame_fifo_wrport_dat_w;
wire [8:0] frame_fifo_rdport_adr;
wire [130:0] frame_fifo_rdport_dat_r;
wire frame_fifo_fifo_in_payload_sof;
wire [127:0] frame_fifo_fifo_in_payload_pixels;
wire frame_fifo_fifo_in_first;
wire frame_fifo_fifo_in_last;
wire frame_fifo_fifo_out_payload_sof;
wire [127:0] frame_fifo_fifo_out_payload_pixels;
wire frame_fifo_fifo_out_first;
wire frame_fifo_fifo_out_last;
reg frame_pix_overflow = 1'd0;
wire frame_pix_overflow_reset;
wire frame_sys_overflow;
wire frame_overflow_reset_i;
wire frame_overflow_reset_o;
reg frame_overflow_reset_toggle_i = 1'd0;
wire frame_overflow_reset_toggle_o;
reg frame_overflow_reset_toggle_o_r = 1'd0;
wire frame_overflow_reset_ack_i;
wire frame_overflow_reset_ack_o;
reg frame_overflow_reset_ack_toggle_i = 1'd0;
wire frame_overflow_reset_ack_toggle_o;
reg frame_overflow_reset_ack_toggle_o_r = 1'd0;
reg frame_overflow_mask = 1'd0;
wire dma_frame_valid;
reg dma_frame_ready = 1'd0;
wire dma_frame_first;
wire dma_frame_last;
wire dma_frame_payload_sof;
wire [127:0] dma_frame_payload_pixels;
reg [28:0] dma_frame_size_storage_full = 29'd0;
wire [24:0] dma_frame_size_storage;
reg dma_frame_size_re = 1'd0;
wire dma_slot_array_irq;
wire [24:0] dma_slot_array_address;
wire [24:0] dma_slot_array_address_reached;
wire dma_slot_array_address_valid;
reg dma_slot_array_address_done = 1'd0;
wire dma_slot_array_slot0_status;
wire dma_slot_array_slot0_pending;
wire dma_slot_array_slot0_trigger;
reg dma_slot_array_slot0_clear = 1'd0;
wire [24:0] dma_slot_array_slot0_address;
wire [24:0] dma_slot_array_slot0_address_reached;
wire dma_slot_array_slot0_address_valid;
wire dma_slot_array_slot0_address_done;
reg [1:0] dma_slot_array_slot0_status_storage_full = 2'd0;
wire [1:0] dma_slot_array_slot0_status_storage;
reg dma_slot_array_slot0_status_re = 1'd0;
wire dma_slot_array_slot0_status_we;
wire [1:0] dma_slot_array_slot0_status_dat_w;
reg [28:0] dma_slot_array_slot0_address_storage_full = 29'd0;
wire [24:0] dma_slot_array_slot0_address_storage;
reg dma_slot_array_slot0_address_re = 1'd0;
wire dma_slot_array_slot0_address_we;
wire [24:0] dma_slot_array_slot0_address_dat_w;
wire dma_slot_array_slot1_status;
wire dma_slot_array_slot1_pending;
wire dma_slot_array_slot1_trigger;
reg dma_slot_array_slot1_clear = 1'd0;
wire [24:0] dma_slot_array_slot1_address;
wire [24:0] dma_slot_array_slot1_address_reached;
wire dma_slot_array_slot1_address_valid;
wire dma_slot_array_slot1_address_done;
reg [1:0] dma_slot_array_slot1_status_storage_full = 2'd0;
wire [1:0] dma_slot_array_slot1_status_storage;
reg dma_slot_array_slot1_status_re = 1'd0;
wire dma_slot_array_slot1_status_we;
wire [1:0] dma_slot_array_slot1_status_dat_w;
reg [28:0] dma_slot_array_slot1_address_storage_full = 29'd0;
wire [24:0] dma_slot_array_slot1_address_storage;
reg dma_slot_array_slot1_address_re = 1'd0;
wire dma_slot_array_slot1_address_we;
wire [24:0] dma_slot_array_slot1_address_dat_w;
wire dma_slot_array_status_re;
wire [1:0] dma_slot_array_status_r;
reg [1:0] dma_slot_array_status_w = 2'd0;
wire dma_slot_array_pending_re;
wire [1:0] dma_slot_array_pending_r;
reg [1:0] dma_slot_array_pending_w = 2'd0;
reg [1:0] dma_slot_array_storage_full = 2'd0;
wire [1:0] dma_slot_array_storage;
reg dma_slot_array_re = 1'd0;
wire dma_slot_array_change_slot;
reg dma_slot_array_current_slot = 1'd0;
reg dma_reset_words = 1'd0;
reg dma_count_word = 1'd0;
wire dma_last_word;
reg [24:0] dma_current_address = 25'd0;
reg [24:0] dma_mwords_remaining = 25'd0;
wire [127:0] dma_memory_word;
reg dma_sink_sink_valid = 1'd0;
wire dma_sink_sink_ready;
wire [24:0] dma_sink_sink_payload_address;
wire [127:0] dma_sink_sink_payload_data;
wire dma_fifo_sink_valid;
wire dma_fifo_sink_ready;
reg dma_fifo_sink_first = 1'd0;
reg dma_fifo_sink_last = 1'd0;
wire [127:0] dma_fifo_sink_payload_data;
wire dma_fifo_source_valid;
wire dma_fifo_source_ready;
wire dma_fifo_source_first;
wire dma_fifo_source_last;
wire [127:0] dma_fifo_source_payload_data;
wire dma_fifo_syncfifo_we;
wire dma_fifo_syncfifo_writable;
wire dma_fifo_syncfifo_re;
wire dma_fifo_syncfifo_readable;
wire [129:0] dma_fifo_syncfifo_din;
wire [129:0] dma_fifo_syncfifo_dout;
reg [4:0] dma_fifo_level = 5'd0;
reg dma_fifo_replace = 1'd0;
reg [3:0] dma_fifo_produce = 4'd0;
reg [3:0] dma_fifo_consume = 4'd0;
reg [3:0] dma_fifo_wrport_adr = 4'd0;
wire [129:0] dma_fifo_wrport_dat_r;
wire dma_fifo_wrport_we;
wire [129:0] dma_fifo_wrport_dat_w;
wire dma_fifo_do_read;
wire [3:0] dma_fifo_rdport_adr;
wire [129:0] dma_fifo_rdport_dat_r;
wire [127:0] dma_fifo_fifo_in_payload_data;
wire dma_fifo_fifo_in_first;
wire dma_fifo_fifo_in_last;
wire [127:0] dma_fifo_fifo_out_payload_data;
wire dma_fifo_fifo_out_first;
wire dma_fifo_fifo_out_last;
wire hdmi_in0_freq_clk0;
wire [31:0] hdmi_in0_freq_status;
wire fmeter_clk;
wire hdmi_in0_freq_period_done;
reg [31:0] hdmi_in0_freq_period_counter = 32'd0;
wire hdmi_in0_freq_ce;
reg [5:0] hdmi_in0_freq_q = 6'd0;
wire [5:0] hdmi_in0_freq_q_next;
reg [5:0] hdmi_in0_freq_q_binary = 6'd0;
reg [5:0] hdmi_in0_freq_q_next_binary = 6'd0;
wire [5:0] hdmi_in0_freq_gray_decoder_i;
reg [5:0] hdmi_in0_freq_gray_decoder_o = 6'd0;
reg [5:0] hdmi_in0_freq_gray_decoder_o_comb = 6'd0;
wire hdmi_in0_freq_sampler_latch;
wire [5:0] hdmi_in0_freq_sampler_i;
reg [31:0] hdmi_in0_freq_sampler_o = 32'd0;
wire [5:0] hdmi_in0_freq_sampler_inc;
reg [31:0] hdmi_in0_freq_sampler_counter = 32'd0;
reg [5:0] hdmi_in0_freq_sampler_i_d = 6'd0;
wire hdmi_out0_dram_port_cmd_valid;
wire hdmi_out0_dram_port_cmd_ready;
wire hdmi_out0_dram_port_cmd_first;
wire hdmi_out0_dram_port_cmd_last;
wire hdmi_out0_dram_port_cmd_payload_we;
wire [24:0] hdmi_out0_dram_port_cmd_payload_adr;
wire hdmi_out0_dram_port_wdata_ready;
reg [127:0] hdmi_out0_dram_port_wdata_payload_data = 128'd0;
reg [15:0] hdmi_out0_dram_port_wdata_payload_we = 16'd0;
wire hdmi_out0_dram_port_rdata_valid;
wire hdmi_out0_dram_port_rdata_ready;
reg hdmi_out0_dram_port_rdata_first = 1'd0;
reg hdmi_out0_dram_port_rdata_last = 1'd0;
wire [127:0] hdmi_out0_dram_port_rdata_payload_data;
reg hdmi_out0_dram_port_litedramport0_cmd_valid = 1'd0;
wire hdmi_out0_dram_port_litedramport0_cmd_ready;
reg hdmi_out0_dram_port_litedramport0_cmd_first = 1'd0;
reg hdmi_out0_dram_port_litedramport0_cmd_last = 1'd0;
reg hdmi_out0_dram_port_litedramport0_cmd_payload_we = 1'd0;
reg [24:0] hdmi_out0_dram_port_litedramport0_cmd_payload_adr = 25'd0;
wire hdmi_out0_dram_port_litedramport0_rdata_valid;
wire hdmi_out0_dram_port_litedramport0_rdata_ready;
wire hdmi_out0_dram_port_litedramport0_rdata_first;
wire hdmi_out0_dram_port_litedramport0_rdata_last;
wire [127:0] hdmi_out0_dram_port_litedramport0_rdata_payload_data;
wire hdmi_out0_dram_port_cmd_fifo_sink_valid;
wire hdmi_out0_dram_port_cmd_fifo_sink_ready;
wire hdmi_out0_dram_port_cmd_fifo_sink_first;
wire hdmi_out0_dram_port_cmd_fifo_sink_last;
wire hdmi_out0_dram_port_cmd_fifo_sink_payload_we;
wire [24:0] hdmi_out0_dram_port_cmd_fifo_sink_payload_adr;
wire hdmi_out0_dram_port_cmd_fifo_source_valid;
wire hdmi_out0_dram_port_cmd_fifo_source_ready;
wire hdmi_out0_dram_port_cmd_fifo_source_first;
wire hdmi_out0_dram_port_cmd_fifo_source_last;
wire hdmi_out0_dram_port_cmd_fifo_source_payload_we;
wire [24:0] hdmi_out0_dram_port_cmd_fifo_source_payload_adr;
wire hdmi_out0_dram_port_cmd_fifo_asyncfifo_we;
wire hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable;
wire hdmi_out0_dram_port_cmd_fifo_asyncfifo_re;
wire hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable;
wire [27:0] hdmi_out0_dram_port_cmd_fifo_asyncfifo_din;
wire [27:0] hdmi_out0_dram_port_cmd_fifo_asyncfifo_dout;
wire hdmi_out0_dram_port_cmd_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter0_q = 3'd0;
wire [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next;
reg [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary = 3'd0;
reg [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary = 3'd0;
wire hdmi_out0_dram_port_cmd_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter1_q = 3'd0;
wire [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next;
reg [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary = 3'd0;
reg [2:0] hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary = 3'd0;
wire [2:0] hdmi_out0_dram_port_cmd_fifo_produce_rdomain;
wire [2:0] hdmi_out0_dram_port_cmd_fifo_consume_wdomain;
wire [1:0] hdmi_out0_dram_port_cmd_fifo_wrport_adr;
wire [27:0] hdmi_out0_dram_port_cmd_fifo_wrport_dat_r;
wire hdmi_out0_dram_port_cmd_fifo_wrport_we;
wire [27:0] hdmi_out0_dram_port_cmd_fifo_wrport_dat_w;
wire [1:0] hdmi_out0_dram_port_cmd_fifo_rdport_adr;
wire [27:0] hdmi_out0_dram_port_cmd_fifo_rdport_dat_r;
wire hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_we;
wire [24:0] hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_adr;
wire hdmi_out0_dram_port_cmd_fifo_fifo_in_first;
wire hdmi_out0_dram_port_cmd_fifo_fifo_in_last;
wire hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_we;
wire [24:0] hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_adr;
wire hdmi_out0_dram_port_cmd_fifo_fifo_out_first;
wire hdmi_out0_dram_port_cmd_fifo_fifo_out_last;
wire hdmi_out0_dram_port_rdata_fifo_sink_valid;
wire hdmi_out0_dram_port_rdata_fifo_sink_ready;
wire hdmi_out0_dram_port_rdata_fifo_sink_first;
wire hdmi_out0_dram_port_rdata_fifo_sink_last;
wire [127:0] hdmi_out0_dram_port_rdata_fifo_sink_payload_data;
wire hdmi_out0_dram_port_rdata_fifo_source_valid;
wire hdmi_out0_dram_port_rdata_fifo_source_ready;
wire hdmi_out0_dram_port_rdata_fifo_source_first;
wire hdmi_out0_dram_port_rdata_fifo_source_last;
wire [127:0] hdmi_out0_dram_port_rdata_fifo_source_payload_data;
wire hdmi_out0_dram_port_rdata_fifo_asyncfifo_we;
wire hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable;
wire hdmi_out0_dram_port_rdata_fifo_asyncfifo_re;
wire hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable;
wire [129:0] hdmi_out0_dram_port_rdata_fifo_asyncfifo_din;
wire [129:0] hdmi_out0_dram_port_rdata_fifo_asyncfifo_dout;
wire hdmi_out0_dram_port_rdata_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter0_q = 5'd0;
wire [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next;
reg [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary = 5'd0;
reg [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary = 5'd0;
wire hdmi_out0_dram_port_rdata_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter1_q = 5'd0;
wire [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next;
reg [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary = 5'd0;
reg [4:0] hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary = 5'd0;
wire [4:0] hdmi_out0_dram_port_rdata_fifo_produce_rdomain;
wire [4:0] hdmi_out0_dram_port_rdata_fifo_consume_wdomain;
wire [3:0] hdmi_out0_dram_port_rdata_fifo_wrport_adr;
wire [129:0] hdmi_out0_dram_port_rdata_fifo_wrport_dat_r;
wire hdmi_out0_dram_port_rdata_fifo_wrport_we;
wire [129:0] hdmi_out0_dram_port_rdata_fifo_wrport_dat_w;
wire [3:0] hdmi_out0_dram_port_rdata_fifo_rdport_adr;
wire [129:0] hdmi_out0_dram_port_rdata_fifo_rdport_dat_r;
wire [127:0] hdmi_out0_dram_port_rdata_fifo_fifo_in_payload_data;
wire hdmi_out0_dram_port_rdata_fifo_fifo_in_first;
wire hdmi_out0_dram_port_rdata_fifo_fifo_in_last;
wire [127:0] hdmi_out0_dram_port_rdata_fifo_fifo_out_payload_data;
wire hdmi_out0_dram_port_rdata_fifo_fifo_out_first;
wire hdmi_out0_dram_port_rdata_fifo_fifo_out_last;
wire hdmi_out0_dram_port_litedramport1_cmd_valid;
reg hdmi_out0_dram_port_litedramport1_cmd_ready = 1'd0;
wire hdmi_out0_dram_port_litedramport1_cmd_payload_we;
wire [27:0] hdmi_out0_dram_port_litedramport1_cmd_payload_adr;
reg hdmi_out0_dram_port_litedramport1_rdata_valid = 1'd0;
wire hdmi_out0_dram_port_litedramport1_rdata_ready;
reg hdmi_out0_dram_port_litedramport1_rdata_first = 1'd0;
reg hdmi_out0_dram_port_litedramport1_rdata_last = 1'd0;
reg [15:0] hdmi_out0_dram_port_litedramport1_rdata_payload_data = 16'd0;
reg hdmi_out0_dram_port_litedramport1_flush = 1'd0;
reg hdmi_out0_dram_port_cmd_buffer_sink_valid = 1'd0;
wire hdmi_out0_dram_port_cmd_buffer_sink_ready;
reg hdmi_out0_dram_port_cmd_buffer_sink_first = 1'd0;
reg hdmi_out0_dram_port_cmd_buffer_sink_last = 1'd0;
reg [7:0] hdmi_out0_dram_port_cmd_buffer_sink_payload_sel = 8'd0;
wire hdmi_out0_dram_port_cmd_buffer_source_valid;
wire hdmi_out0_dram_port_cmd_buffer_source_ready;
wire hdmi_out0_dram_port_cmd_buffer_source_first;
wire hdmi_out0_dram_port_cmd_buffer_source_last;
wire [7:0] hdmi_out0_dram_port_cmd_buffer_source_payload_sel;
wire hdmi_out0_dram_port_cmd_buffer_syncfifo_we;
wire hdmi_out0_dram_port_cmd_buffer_syncfifo_writable;
wire hdmi_out0_dram_port_cmd_buffer_syncfifo_re;
wire hdmi_out0_dram_port_cmd_buffer_syncfifo_readable;
wire [9:0] hdmi_out0_dram_port_cmd_buffer_syncfifo_din;
wire [9:0] hdmi_out0_dram_port_cmd_buffer_syncfifo_dout;
reg [2:0] hdmi_out0_dram_port_cmd_buffer_level = 3'd0;
reg hdmi_out0_dram_port_cmd_buffer_replace = 1'd0;
reg [1:0] hdmi_out0_dram_port_cmd_buffer_produce = 2'd0;
reg [1:0] hdmi_out0_dram_port_cmd_buffer_consume = 2'd0;
reg [1:0] hdmi_out0_dram_port_cmd_buffer_wrport_adr = 2'd0;
wire [9:0] hdmi_out0_dram_port_cmd_buffer_wrport_dat_r;
wire hdmi_out0_dram_port_cmd_buffer_wrport_we;
wire [9:0] hdmi_out0_dram_port_cmd_buffer_wrport_dat_w;
wire hdmi_out0_dram_port_cmd_buffer_do_read;
wire [1:0] hdmi_out0_dram_port_cmd_buffer_rdport_adr;
wire [9:0] hdmi_out0_dram_port_cmd_buffer_rdport_dat_r;
wire [7:0] hdmi_out0_dram_port_cmd_buffer_fifo_in_payload_sel;
wire hdmi_out0_dram_port_cmd_buffer_fifo_in_first;
wire hdmi_out0_dram_port_cmd_buffer_fifo_in_last;
wire [7:0] hdmi_out0_dram_port_cmd_buffer_fifo_out_payload_sel;
wire hdmi_out0_dram_port_cmd_buffer_fifo_out_first;
wire hdmi_out0_dram_port_cmd_buffer_fifo_out_last;
reg [2:0] hdmi_out0_dram_port_counter = 3'd0;
reg hdmi_out0_dram_port_counter_ce = 1'd0;
wire hdmi_out0_dram_port_rdata_buffer_sink_valid;
wire hdmi_out0_dram_port_rdata_buffer_sink_ready;
wire hdmi_out0_dram_port_rdata_buffer_sink_first;
wire hdmi_out0_dram_port_rdata_buffer_sink_last;
wire [127:0] hdmi_out0_dram_port_rdata_buffer_sink_payload_data;
wire hdmi_out0_dram_port_rdata_buffer_source_valid;
wire hdmi_out0_dram_port_rdata_buffer_source_ready;
wire hdmi_out0_dram_port_rdata_buffer_source_first;
wire hdmi_out0_dram_port_rdata_buffer_source_last;
reg [127:0] hdmi_out0_dram_port_rdata_buffer_source_payload_data = 128'd0;
wire hdmi_out0_dram_port_rdata_buffer_pipe_ce;
wire hdmi_out0_dram_port_rdata_buffer_busy;
reg hdmi_out0_dram_port_rdata_buffer_valid_n = 1'd0;
reg hdmi_out0_dram_port_rdata_buffer_first_n = 1'd0;
reg hdmi_out0_dram_port_rdata_buffer_last_n = 1'd0;
wire hdmi_out0_dram_port_rdata_converter_sink_valid;
wire hdmi_out0_dram_port_rdata_converter_sink_ready;
wire hdmi_out0_dram_port_rdata_converter_sink_first;
wire hdmi_out0_dram_port_rdata_converter_sink_last;
wire [127:0] hdmi_out0_dram_port_rdata_converter_sink_payload_data;
wire hdmi_out0_dram_port_rdata_converter_source_valid;
reg hdmi_out0_dram_port_rdata_converter_source_ready = 1'd0;
wire hdmi_out0_dram_port_rdata_converter_source_first;
wire hdmi_out0_dram_port_rdata_converter_source_last;
wire [15:0] hdmi_out0_dram_port_rdata_converter_source_payload_data;
wire hdmi_out0_dram_port_rdata_converter_converter_sink_valid;
wire hdmi_out0_dram_port_rdata_converter_converter_sink_ready;
wire hdmi_out0_dram_port_rdata_converter_converter_sink_first;
wire hdmi_out0_dram_port_rdata_converter_converter_sink_last;
reg [127:0] hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data = 128'd0;
wire hdmi_out0_dram_port_rdata_converter_converter_source_valid;
wire hdmi_out0_dram_port_rdata_converter_converter_source_ready;
wire hdmi_out0_dram_port_rdata_converter_converter_source_first;
wire hdmi_out0_dram_port_rdata_converter_converter_source_last;
reg [15:0] hdmi_out0_dram_port_rdata_converter_converter_source_payload_data = 16'd0;
wire hdmi_out0_dram_port_rdata_converter_converter_source_payload_valid_token_count;
reg [2:0] hdmi_out0_dram_port_rdata_converter_converter_mux = 3'd0;
wire hdmi_out0_dram_port_rdata_converter_converter_first;
wire hdmi_out0_dram_port_rdata_converter_converter_last;
wire hdmi_out0_dram_port_rdata_converter_source_source_valid;
wire hdmi_out0_dram_port_rdata_converter_source_source_ready;
wire hdmi_out0_dram_port_rdata_converter_source_source_first;
wire hdmi_out0_dram_port_rdata_converter_source_source_last;
wire [15:0] hdmi_out0_dram_port_rdata_converter_source_source_payload_data;
reg [7:0] hdmi_out0_dram_port_rdata_chunk = 8'd1;
wire hdmi_out0_dram_port_rdata_chunk_valid;
wire hdmi_out0_core_source_source_valid;
wire hdmi_out0_core_source_source_ready;
wire [15:0] hdmi_out0_core_source_source_payload_data;
wire hdmi_out0_core_source_source_param_hsync;
wire hdmi_out0_core_source_source_param_vsync;
wire hdmi_out0_core_source_source_param_de;
reg hdmi_out0_core_underflow_enable_storage_full = 1'd0;
wire hdmi_out0_core_underflow_enable_storage;
reg hdmi_out0_core_underflow_enable_re = 1'd0;
wire hdmi_out0_core_underflow_update_underflow_update_re;
wire hdmi_out0_core_underflow_update_underflow_update_r;
reg hdmi_out0_core_underflow_update_underflow_update_w = 1'd0;
reg [31:0] hdmi_out0_core_underflow_counter_status = 32'd0;
wire hdmi_out0_core_initiator_source_source_valid;
wire hdmi_out0_core_initiator_source_source_ready;
wire hdmi_out0_core_initiator_source_source_first;
wire hdmi_out0_core_initiator_source_source_last;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_hres;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_hsync_start;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_hsync_end;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_hscan;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_vres;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_vsync_start;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_vsync_end;
wire [11:0] hdmi_out0_core_initiator_source_source_payload_vscan;
wire [31:0] hdmi_out0_core_initiator_source_source_payload_base;
wire [31:0] hdmi_out0_core_initiator_source_source_payload_length;
wire hdmi_out0_core_initiator_cdc_sink_valid;
wire hdmi_out0_core_initiator_cdc_sink_ready;
reg hdmi_out0_core_initiator_cdc_sink_first = 1'd0;
reg hdmi_out0_core_initiator_cdc_sink_last = 1'd0;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_hres;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_hsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_hsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_hscan;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_vres;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_vsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_vsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_sink_payload_vscan;
wire [31:0] hdmi_out0_core_initiator_cdc_sink_payload_base;
wire [31:0] hdmi_out0_core_initiator_cdc_sink_payload_length;
wire hdmi_out0_core_initiator_cdc_source_valid;
wire hdmi_out0_core_initiator_cdc_source_ready;
wire hdmi_out0_core_initiator_cdc_source_first;
wire hdmi_out0_core_initiator_cdc_source_last;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_hres;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_hsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_hsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_hscan;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_vres;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_vsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_vsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_source_payload_vscan;
wire [31:0] hdmi_out0_core_initiator_cdc_source_payload_base;
wire [31:0] hdmi_out0_core_initiator_cdc_source_payload_length;
wire hdmi_out0_core_initiator_cdc_asyncfifo_we;
wire hdmi_out0_core_initiator_cdc_asyncfifo_writable;
wire hdmi_out0_core_initiator_cdc_asyncfifo_re;
wire hdmi_out0_core_initiator_cdc_asyncfifo_readable;
wire [161:0] hdmi_out0_core_initiator_cdc_asyncfifo_din;
wire [161:0] hdmi_out0_core_initiator_cdc_asyncfifo_dout;
wire hdmi_out0_core_initiator_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [1:0] hdmi_out0_core_initiator_cdc_graycounter0_q = 2'd0;
wire [1:0] hdmi_out0_core_initiator_cdc_graycounter0_q_next;
reg [1:0] hdmi_out0_core_initiator_cdc_graycounter0_q_binary = 2'd0;
reg [1:0] hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary = 2'd0;
wire hdmi_out0_core_initiator_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [1:0] hdmi_out0_core_initiator_cdc_graycounter1_q = 2'd0;
wire [1:0] hdmi_out0_core_initiator_cdc_graycounter1_q_next;
reg [1:0] hdmi_out0_core_initiator_cdc_graycounter1_q_binary = 2'd0;
reg [1:0] hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary = 2'd0;
wire [1:0] hdmi_out0_core_initiator_cdc_produce_rdomain;
wire [1:0] hdmi_out0_core_initiator_cdc_consume_wdomain;
wire hdmi_out0_core_initiator_cdc_wrport_adr;
wire [161:0] hdmi_out0_core_initiator_cdc_wrport_dat_r;
wire hdmi_out0_core_initiator_cdc_wrport_we;
wire [161:0] hdmi_out0_core_initiator_cdc_wrport_dat_w;
wire hdmi_out0_core_initiator_cdc_rdport_adr;
wire [161:0] hdmi_out0_core_initiator_cdc_rdport_dat_r;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_hres;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_vres;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan;
wire [31:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_base;
wire [31:0] hdmi_out0_core_initiator_cdc_fifo_in_payload_length;
wire hdmi_out0_core_initiator_cdc_fifo_in_first;
wire hdmi_out0_core_initiator_cdc_fifo_in_last;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_hres;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_vres;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end;
wire [11:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan;
wire [31:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_base;
wire [31:0] hdmi_out0_core_initiator_cdc_fifo_out_payload_length;
wire hdmi_out0_core_initiator_cdc_fifo_out_first;
wire hdmi_out0_core_initiator_cdc_fifo_out_last;
reg hdmi_out0_core_initiator_enable_storage_full = 1'd0;
wire hdmi_out0_core_initiator_enable_storage;
reg hdmi_out0_core_initiator_enable_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage0_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage0_storage;
reg hdmi_out0_core_initiator_csrstorage0_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage1_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage1_storage;
reg hdmi_out0_core_initiator_csrstorage1_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage2_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage2_storage;
reg hdmi_out0_core_initiator_csrstorage2_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage3_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage3_storage;
reg hdmi_out0_core_initiator_csrstorage3_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage4_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage4_storage;
reg hdmi_out0_core_initiator_csrstorage4_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage5_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage5_storage;
reg hdmi_out0_core_initiator_csrstorage5_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage6_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage6_storage;
reg hdmi_out0_core_initiator_csrstorage6_re = 1'd0;
reg [11:0] hdmi_out0_core_initiator_csrstorage7_storage_full = 12'd0;
wire [11:0] hdmi_out0_core_initiator_csrstorage7_storage;
reg hdmi_out0_core_initiator_csrstorage7_re = 1'd0;
reg [31:0] hdmi_out0_core_initiator_csrstorage8_storage_full = 32'd0;
wire [31:0] hdmi_out0_core_initiator_csrstorage8_storage;
reg hdmi_out0_core_initiator_csrstorage8_re = 1'd0;
reg [31:0] hdmi_out0_core_initiator_csrstorage9_storage_full = 32'd0;
wire [31:0] hdmi_out0_core_initiator_csrstorage9_storage;
reg hdmi_out0_core_initiator_csrstorage9_re = 1'd0;
wire hdmi_out0_core_timinggenerator_sink_valid;
wire hdmi_out0_core_timinggenerator_sink_ready;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_hres;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_hsync_start;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_hsync_end;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_hscan;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_vres;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_vsync_start;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_vsync_end;
wire [11:0] hdmi_out0_core_timinggenerator_sink_payload_vscan;
reg hdmi_out0_core_timinggenerator_source_valid = 1'd0;
reg hdmi_out0_core_timinggenerator_source_ready = 1'd0;
reg hdmi_out0_core_timinggenerator_source_last = 1'd0;
reg hdmi_out0_core_timinggenerator_source_payload_hsync = 1'd0;
reg hdmi_out0_core_timinggenerator_source_payload_vsync = 1'd0;
reg hdmi_out0_core_timinggenerator_source_payload_de = 1'd0;
reg hdmi_out0_core_timinggenerator_hactive = 1'd0;
reg hdmi_out0_core_timinggenerator_vactive = 1'd0;
reg hdmi_out0_core_timinggenerator_active = 1'd0;
reg [11:0] hdmi_out0_core_timinggenerator_hcounter = 12'd0;
reg [11:0] hdmi_out0_core_timinggenerator_vcounter = 12'd0;
wire hdmi_out0_core_dmareader_sink_valid;
reg hdmi_out0_core_dmareader_sink_ready = 1'd0;
wire [31:0] hdmi_out0_core_dmareader_sink_payload_base;
wire [31:0] hdmi_out0_core_dmareader_sink_payload_length;
wire hdmi_out0_core_dmareader_source_valid;
reg hdmi_out0_core_dmareader_source_ready = 1'd0;
wire hdmi_out0_core_dmareader_source_first;
wire hdmi_out0_core_dmareader_source_last;
wire [15:0] hdmi_out0_core_dmareader_source_payload_data;
reg hdmi_out0_core_dmareader_sink_sink_valid = 1'd0;
wire hdmi_out0_core_dmareader_sink_sink_ready;
wire [27:0] hdmi_out0_core_dmareader_sink_sink_payload_address;
wire hdmi_out0_core_dmareader_source_source_valid;
wire hdmi_out0_core_dmareader_source_source_ready;
wire hdmi_out0_core_dmareader_source_source_first;
wire hdmi_out0_core_dmareader_source_source_last;
wire [15:0] hdmi_out0_core_dmareader_source_source_payload_data;
wire hdmi_out0_core_dmareader_request_enable;
wire hdmi_out0_core_dmareader_request_issued;
wire hdmi_out0_core_dmareader_data_dequeued;
reg [12:0] hdmi_out0_core_dmareader_rsv_level = 13'd0;
wire hdmi_out0_core_dmareader_fifo_sink_valid;
wire hdmi_out0_core_dmareader_fifo_sink_ready;
wire hdmi_out0_core_dmareader_fifo_sink_first;
wire hdmi_out0_core_dmareader_fifo_sink_last;
wire [15:0] hdmi_out0_core_dmareader_fifo_sink_payload_data;
wire hdmi_out0_core_dmareader_fifo_source_valid;
wire hdmi_out0_core_dmareader_fifo_source_ready;
wire hdmi_out0_core_dmareader_fifo_source_first;
wire hdmi_out0_core_dmareader_fifo_source_last;
wire [15:0] hdmi_out0_core_dmareader_fifo_source_payload_data;
wire hdmi_out0_core_dmareader_fifo_re;
reg hdmi_out0_core_dmareader_fifo_readable = 1'd0;
wire hdmi_out0_core_dmareader_fifo_syncfifo_we;
wire hdmi_out0_core_dmareader_fifo_syncfifo_writable;
wire hdmi_out0_core_dmareader_fifo_syncfifo_re;
wire hdmi_out0_core_dmareader_fifo_syncfifo_readable;
wire [17:0] hdmi_out0_core_dmareader_fifo_syncfifo_din;
wire [17:0] hdmi_out0_core_dmareader_fifo_syncfifo_dout;
reg [12:0] hdmi_out0_core_dmareader_fifo_level0 = 13'd0;
reg hdmi_out0_core_dmareader_fifo_replace = 1'd0;
reg [11:0] hdmi_out0_core_dmareader_fifo_produce = 12'd0;
reg [11:0] hdmi_out0_core_dmareader_fifo_consume = 12'd0;
reg [11:0] hdmi_out0_core_dmareader_fifo_wrport_adr = 12'd0;
wire [17:0] hdmi_out0_core_dmareader_fifo_wrport_dat_r;
wire hdmi_out0_core_dmareader_fifo_wrport_we;
wire [17:0] hdmi_out0_core_dmareader_fifo_wrport_dat_w;
wire hdmi_out0_core_dmareader_fifo_do_read;
wire [11:0] hdmi_out0_core_dmareader_fifo_rdport_adr;
wire [17:0] hdmi_out0_core_dmareader_fifo_rdport_dat_r;
wire hdmi_out0_core_dmareader_fifo_rdport_re;
wire [12:0] hdmi_out0_core_dmareader_fifo_level1;
wire [15:0] hdmi_out0_core_dmareader_fifo_fifo_in_payload_data;
wire hdmi_out0_core_dmareader_fifo_fifo_in_first;
wire hdmi_out0_core_dmareader_fifo_fifo_in_last;
wire [15:0] hdmi_out0_core_dmareader_fifo_fifo_out_payload_data;
wire hdmi_out0_core_dmareader_fifo_fifo_out_first;
wire hdmi_out0_core_dmareader_fifo_fifo_out_last;
wire [27:0] hdmi_out0_core_dmareader_base;
wire [27:0] hdmi_out0_core_dmareader_length;
reg [27:0] hdmi_out0_core_dmareader_offset = 28'd0;
wire hdmi_out0_core_underflow_enable;
wire hdmi_out0_core_underflow_update;
reg [31:0] hdmi_out0_core_underflow_counter = 32'd0;
wire hdmi_out0_core_i;
wire hdmi_out0_core_o;
reg hdmi_out0_core_toggle_i = 1'd0;
wire hdmi_out0_core_toggle_o;
reg hdmi_out0_core_toggle_o_r = 1'd0;
wire hdmi_out0_driver_sink_sink_valid;
wire hdmi_out0_driver_sink_sink_ready;
wire hdmi_out0_driver_sink_sink_first;
wire hdmi_out0_driver_sink_sink_last;
wire [7:0] hdmi_out0_driver_sink_sink_payload_r;
wire [7:0] hdmi_out0_driver_sink_sink_payload_g;
wire [7:0] hdmi_out0_driver_sink_sink_payload_b;
wire hdmi_out0_driver_sink_sink_param_hsync;
wire hdmi_out0_driver_sink_sink_param_vsync;
wire hdmi_out0_driver_sink_sink_param_de;
wire hdmi_out0_pix_clk;
wire hdmi_out0_pix_rst;
wire hdmi_out0_pix5x_clk;
reg hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full = 1'd0;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage;
reg hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_re = 1'd0;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_read_r;
reg hdmi_out0_driver_s7hdmioutclocking_mmcm_read_w = 1'd0;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_write_r;
reg hdmi_out0_driver_s7hdmioutclocking_mmcm_write_w = 1'd0;
reg hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status = 1'd0;
reg [6:0] hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full = 7'd0;
wire [6:0] hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage;
reg hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_re = 1'd0;
reg [15:0] hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full = 16'd0;
wire [15:0] hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage;
reg hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_re = 1'd0;
wire [15:0] hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_locked;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_fb;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_clk0;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_clk1;
wire hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy;
wire [9:0] hdmi_out0_driver_s7hdmioutclocking_data0;
wire [9:0] hdmi_out0_driver_s7hdmioutclocking_data1;
reg hdmi_out0_driver_s7hdmioutclocking_ce = 1'd0;
wire [1:0] hdmi_out0_driver_s7hdmioutclocking_shift;
wire hdmi_out0_driver_s7hdmioutclocking_pad_se;
reg [9:0] hdmi_out0_driver_s7hdmioutclocking = 10'd31;
wire hdmi_out0_driver_hdmi_phy_sink_valid;
wire hdmi_out0_driver_hdmi_phy_sink_ready;
wire hdmi_out0_driver_hdmi_phy_sink_first;
wire hdmi_out0_driver_hdmi_phy_sink_last;
wire [7:0] hdmi_out0_driver_hdmi_phy_sink_payload_r;
wire [7:0] hdmi_out0_driver_hdmi_phy_sink_payload_g;
wire [7:0] hdmi_out0_driver_hdmi_phy_sink_payload_b;
wire hdmi_out0_driver_hdmi_phy_sink_param_hsync;
wire hdmi_out0_driver_hdmi_phy_sink_param_vsync;
wire hdmi_out0_driver_hdmi_phy_sink_param_de;
wire [7:0] hdmi_out0_driver_hdmi_phy_es0_d0;
wire [1:0] hdmi_out0_driver_hdmi_phy_es0_c;
wire hdmi_out0_driver_hdmi_phy_es0_de;
reg [9:0] hdmi_out0_driver_hdmi_phy_es0_out = 10'd0;
reg [7:0] hdmi_out0_driver_hdmi_phy_es0_d1 = 8'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es0_n1d = 4'd0;
reg [8:0] hdmi_out0_driver_hdmi_phy_es0_q_m = 9'd0;
wire hdmi_out0_driver_hdmi_phy_es0_q_m8_n;
reg [8:0] hdmi_out0_driver_hdmi_phy_es0_q_m_r = 9'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es0_n0q_m = 4'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es0_n1q_m = 4'd0;
reg signed [5:0] hdmi_out0_driver_hdmi_phy_es0_cnt = 6'sd64;
reg [1:0] hdmi_out0_driver_hdmi_phy_es0_new_c0 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es0_new_de0 = 1'd0;
reg [1:0] hdmi_out0_driver_hdmi_phy_es0_new_c1 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es0_new_de1 = 1'd0;
reg [1:0] hdmi_out0_driver_hdmi_phy_es0_new_c2 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es0_new_de2 = 1'd0;
wire [9:0] hdmi_out0_driver_hdmi_phy_es0_data;
reg hdmi_out0_driver_hdmi_phy_es0_ce = 1'd0;
wire [1:0] hdmi_out0_driver_hdmi_phy_es0_shift;
wire hdmi_out0_driver_hdmi_phy_es0_pad_se;
wire [7:0] hdmi_out0_driver_hdmi_phy_es1_d0;
wire [1:0] hdmi_out0_driver_hdmi_phy_es1_c;
wire hdmi_out0_driver_hdmi_phy_es1_de;
reg [9:0] hdmi_out0_driver_hdmi_phy_es1_out = 10'd0;
reg [7:0] hdmi_out0_driver_hdmi_phy_es1_d1 = 8'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es1_n1d = 4'd0;
reg [8:0] hdmi_out0_driver_hdmi_phy_es1_q_m = 9'd0;
wire hdmi_out0_driver_hdmi_phy_es1_q_m8_n;
reg [8:0] hdmi_out0_driver_hdmi_phy_es1_q_m_r = 9'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es1_n0q_m = 4'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es1_n1q_m = 4'd0;
reg signed [5:0] hdmi_out0_driver_hdmi_phy_es1_cnt = 6'sd64;
reg [1:0] hdmi_out0_driver_hdmi_phy_es1_new_c0 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es1_new_de0 = 1'd0;
reg [1:0] hdmi_out0_driver_hdmi_phy_es1_new_c1 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es1_new_de1 = 1'd0;
reg [1:0] hdmi_out0_driver_hdmi_phy_es1_new_c2 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es1_new_de2 = 1'd0;
wire [9:0] hdmi_out0_driver_hdmi_phy_es1_data;
reg hdmi_out0_driver_hdmi_phy_es1_ce = 1'd0;
wire [1:0] hdmi_out0_driver_hdmi_phy_es1_shift;
wire hdmi_out0_driver_hdmi_phy_es1_pad_se;
wire [7:0] hdmi_out0_driver_hdmi_phy_es2_d0;
wire [1:0] hdmi_out0_driver_hdmi_phy_es2_c;
wire hdmi_out0_driver_hdmi_phy_es2_de;
reg [9:0] hdmi_out0_driver_hdmi_phy_es2_out = 10'd0;
reg [7:0] hdmi_out0_driver_hdmi_phy_es2_d1 = 8'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es2_n1d = 4'd0;
reg [8:0] hdmi_out0_driver_hdmi_phy_es2_q_m = 9'd0;
wire hdmi_out0_driver_hdmi_phy_es2_q_m8_n;
reg [8:0] hdmi_out0_driver_hdmi_phy_es2_q_m_r = 9'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es2_n0q_m = 4'd0;
reg [3:0] hdmi_out0_driver_hdmi_phy_es2_n1q_m = 4'd0;
reg signed [5:0] hdmi_out0_driver_hdmi_phy_es2_cnt = 6'sd64;
reg [1:0] hdmi_out0_driver_hdmi_phy_es2_new_c0 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es2_new_de0 = 1'd0;
reg [1:0] hdmi_out0_driver_hdmi_phy_es2_new_c1 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es2_new_de1 = 1'd0;
reg [1:0] hdmi_out0_driver_hdmi_phy_es2_new_c2 = 2'd0;
reg hdmi_out0_driver_hdmi_phy_es2_new_de2 = 1'd0;
wire [9:0] hdmi_out0_driver_hdmi_phy_es2_data;
reg hdmi_out0_driver_hdmi_phy_es2_ce = 1'd0;
wire [1:0] hdmi_out0_driver_hdmi_phy_es2_shift;
wire hdmi_out0_driver_hdmi_phy_es2_pad_se;
wire hdmi_out0_resetinserter_sink_sink_valid;
reg hdmi_out0_resetinserter_sink_sink_ready = 1'd0;
wire [7:0] hdmi_out0_resetinserter_sink_sink_payload_y;
wire [7:0] hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
wire hdmi_out0_resetinserter_source_source_valid;
wire hdmi_out0_resetinserter_source_source_ready;
reg hdmi_out0_resetinserter_source_source_first = 1'd0;
reg hdmi_out0_resetinserter_source_source_last = 1'd0;
wire [7:0] hdmi_out0_resetinserter_source_source_payload_y;
wire [7:0] hdmi_out0_resetinserter_source_source_payload_cb;
wire [7:0] hdmi_out0_resetinserter_source_source_payload_cr;
reg hdmi_out0_resetinserter_y_fifo_sink_valid = 1'd0;
wire hdmi_out0_resetinserter_y_fifo_sink_ready;
reg hdmi_out0_resetinserter_y_fifo_sink_first = 1'd0;
reg hdmi_out0_resetinserter_y_fifo_sink_last = 1'd0;
reg [7:0] hdmi_out0_resetinserter_y_fifo_sink_payload_data = 8'd0;
wire hdmi_out0_resetinserter_y_fifo_source_valid;
wire hdmi_out0_resetinserter_y_fifo_source_ready;
wire hdmi_out0_resetinserter_y_fifo_source_first;
wire hdmi_out0_resetinserter_y_fifo_source_last;
wire [7:0] hdmi_out0_resetinserter_y_fifo_source_payload_data;
wire hdmi_out0_resetinserter_y_fifo_syncfifo_we;
wire hdmi_out0_resetinserter_y_fifo_syncfifo_writable;
wire hdmi_out0_resetinserter_y_fifo_syncfifo_re;
wire hdmi_out0_resetinserter_y_fifo_syncfifo_readable;
wire [9:0] hdmi_out0_resetinserter_y_fifo_syncfifo_din;
wire [9:0] hdmi_out0_resetinserter_y_fifo_syncfifo_dout;
reg [2:0] hdmi_out0_resetinserter_y_fifo_level = 3'd0;
reg hdmi_out0_resetinserter_y_fifo_replace = 1'd0;
reg [1:0] hdmi_out0_resetinserter_y_fifo_produce = 2'd0;
reg [1:0] hdmi_out0_resetinserter_y_fifo_consume = 2'd0;
reg [1:0] hdmi_out0_resetinserter_y_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi_out0_resetinserter_y_fifo_wrport_dat_r;
wire hdmi_out0_resetinserter_y_fifo_wrport_we;
wire [9:0] hdmi_out0_resetinserter_y_fifo_wrport_dat_w;
wire hdmi_out0_resetinserter_y_fifo_do_read;
wire [1:0] hdmi_out0_resetinserter_y_fifo_rdport_adr;
wire [9:0] hdmi_out0_resetinserter_y_fifo_rdport_dat_r;
wire [7:0] hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data;
wire hdmi_out0_resetinserter_y_fifo_fifo_in_first;
wire hdmi_out0_resetinserter_y_fifo_fifo_in_last;
wire [7:0] hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data;
wire hdmi_out0_resetinserter_y_fifo_fifo_out_first;
wire hdmi_out0_resetinserter_y_fifo_fifo_out_last;
reg hdmi_out0_resetinserter_cb_fifo_sink_valid = 1'd0;
wire hdmi_out0_resetinserter_cb_fifo_sink_ready;
reg hdmi_out0_resetinserter_cb_fifo_sink_first = 1'd0;
reg hdmi_out0_resetinserter_cb_fifo_sink_last = 1'd0;
reg [7:0] hdmi_out0_resetinserter_cb_fifo_sink_payload_data = 8'd0;
wire hdmi_out0_resetinserter_cb_fifo_source_valid;
wire hdmi_out0_resetinserter_cb_fifo_source_ready;
wire hdmi_out0_resetinserter_cb_fifo_source_first;
wire hdmi_out0_resetinserter_cb_fifo_source_last;
wire [7:0] hdmi_out0_resetinserter_cb_fifo_source_payload_data;
wire hdmi_out0_resetinserter_cb_fifo_syncfifo_we;
wire hdmi_out0_resetinserter_cb_fifo_syncfifo_writable;
wire hdmi_out0_resetinserter_cb_fifo_syncfifo_re;
wire hdmi_out0_resetinserter_cb_fifo_syncfifo_readable;
wire [9:0] hdmi_out0_resetinserter_cb_fifo_syncfifo_din;
wire [9:0] hdmi_out0_resetinserter_cb_fifo_syncfifo_dout;
reg [2:0] hdmi_out0_resetinserter_cb_fifo_level = 3'd0;
reg hdmi_out0_resetinserter_cb_fifo_replace = 1'd0;
reg [1:0] hdmi_out0_resetinserter_cb_fifo_produce = 2'd0;
reg [1:0] hdmi_out0_resetinserter_cb_fifo_consume = 2'd0;
reg [1:0] hdmi_out0_resetinserter_cb_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi_out0_resetinserter_cb_fifo_wrport_dat_r;
wire hdmi_out0_resetinserter_cb_fifo_wrport_we;
wire [9:0] hdmi_out0_resetinserter_cb_fifo_wrport_dat_w;
wire hdmi_out0_resetinserter_cb_fifo_do_read;
wire [1:0] hdmi_out0_resetinserter_cb_fifo_rdport_adr;
wire [9:0] hdmi_out0_resetinserter_cb_fifo_rdport_dat_r;
wire [7:0] hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data;
wire hdmi_out0_resetinserter_cb_fifo_fifo_in_first;
wire hdmi_out0_resetinserter_cb_fifo_fifo_in_last;
wire [7:0] hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data;
wire hdmi_out0_resetinserter_cb_fifo_fifo_out_first;
wire hdmi_out0_resetinserter_cb_fifo_fifo_out_last;
reg hdmi_out0_resetinserter_cr_fifo_sink_valid = 1'd0;
wire hdmi_out0_resetinserter_cr_fifo_sink_ready;
reg hdmi_out0_resetinserter_cr_fifo_sink_first = 1'd0;
reg hdmi_out0_resetinserter_cr_fifo_sink_last = 1'd0;
reg [7:0] hdmi_out0_resetinserter_cr_fifo_sink_payload_data = 8'd0;
wire hdmi_out0_resetinserter_cr_fifo_source_valid;
wire hdmi_out0_resetinserter_cr_fifo_source_ready;
wire hdmi_out0_resetinserter_cr_fifo_source_first;
wire hdmi_out0_resetinserter_cr_fifo_source_last;
wire [7:0] hdmi_out0_resetinserter_cr_fifo_source_payload_data;
wire hdmi_out0_resetinserter_cr_fifo_syncfifo_we;
wire hdmi_out0_resetinserter_cr_fifo_syncfifo_writable;
wire hdmi_out0_resetinserter_cr_fifo_syncfifo_re;
wire hdmi_out0_resetinserter_cr_fifo_syncfifo_readable;
wire [9:0] hdmi_out0_resetinserter_cr_fifo_syncfifo_din;
wire [9:0] hdmi_out0_resetinserter_cr_fifo_syncfifo_dout;
reg [2:0] hdmi_out0_resetinserter_cr_fifo_level = 3'd0;
reg hdmi_out0_resetinserter_cr_fifo_replace = 1'd0;
reg [1:0] hdmi_out0_resetinserter_cr_fifo_produce = 2'd0;
reg [1:0] hdmi_out0_resetinserter_cr_fifo_consume = 2'd0;
reg [1:0] hdmi_out0_resetinserter_cr_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi_out0_resetinserter_cr_fifo_wrport_dat_r;
wire hdmi_out0_resetinserter_cr_fifo_wrport_we;
wire [9:0] hdmi_out0_resetinserter_cr_fifo_wrport_dat_w;
wire hdmi_out0_resetinserter_cr_fifo_do_read;
wire [1:0] hdmi_out0_resetinserter_cr_fifo_rdport_adr;
wire [9:0] hdmi_out0_resetinserter_cr_fifo_rdport_dat_r;
wire [7:0] hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data;
wire hdmi_out0_resetinserter_cr_fifo_fifo_in_first;
wire hdmi_out0_resetinserter_cr_fifo_fifo_in_last;
wire [7:0] hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data;
wire hdmi_out0_resetinserter_cr_fifo_fifo_out_first;
wire hdmi_out0_resetinserter_cr_fifo_fifo_out_last;
reg hdmi_out0_resetinserter_parity_in = 1'd0;
reg hdmi_out0_resetinserter_parity_out = 1'd0;
wire hdmi_out0_resetinserter_reset;
wire hdmi_out0_sink_valid;
wire hdmi_out0_sink_ready;
wire hdmi_out0_sink_first;
wire hdmi_out0_sink_last;
wire [7:0] hdmi_out0_sink_payload_y;
wire [7:0] hdmi_out0_sink_payload_cb;
wire [7:0] hdmi_out0_sink_payload_cr;
wire hdmi_out0_source_valid;
wire hdmi_out0_source_ready;
wire hdmi_out0_source_first;
wire hdmi_out0_source_last;
wire [7:0] hdmi_out0_source_payload_r;
wire [7:0] hdmi_out0_source_payload_g;
wire [7:0] hdmi_out0_source_payload_b;
wire [7:0] hdmi_out0_sink_y;
wire [7:0] hdmi_out0_sink_cb;
wire [7:0] hdmi_out0_sink_cr;
reg [7:0] hdmi_out0_source_r = 8'd0;
reg [7:0] hdmi_out0_source_g = 8'd0;
reg [7:0] hdmi_out0_source_b = 8'd0;
reg [7:0] hdmi_out0_record0_ycbcr_n_y = 8'd0;
reg [7:0] hdmi_out0_record0_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi_out0_record0_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi_out0_record1_ycbcr_n_y = 8'd0;
reg [7:0] hdmi_out0_record1_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi_out0_record1_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi_out0_record2_ycbcr_n_y = 8'd0;
reg [7:0] hdmi_out0_record2_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi_out0_record2_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi_out0_record3_ycbcr_n_y = 8'd0;
reg [7:0] hdmi_out0_record3_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi_out0_record3_ycbcr_n_cr = 8'd0;
reg signed [8:0] hdmi_out0_cb_minus_coffset = 9'sd512;
reg signed [8:0] hdmi_out0_cr_minus_coffset = 9'sd512;
reg signed [8:0] hdmi_out0_y_minus_yoffset = 9'sd512;
reg signed [19:0] hdmi_out0_cr_minus_coffset_mult_acoef = 20'sd1048576;
reg signed [19:0] hdmi_out0_cb_minus_coffset_mult_bcoef = 20'sd1048576;
reg signed [19:0] hdmi_out0_cr_minus_coffset_mult_ccoef = 20'sd1048576;
reg signed [19:0] hdmi_out0_cb_minus_coffset_mult_dcoef = 20'sd1048576;
reg signed [11:0] hdmi_out0_r = 12'sd4096;
reg signed [11:0] hdmi_out0_g = 12'sd4096;
reg signed [11:0] hdmi_out0_b = 12'sd4096;
wire hdmi_out0_ce;
wire hdmi_out0_pipe_ce;
wire hdmi_out0_busy;
reg hdmi_out0_valid_n0 = 1'd0;
reg hdmi_out0_valid_n1 = 1'd0;
reg hdmi_out0_valid_n2 = 1'd0;
reg hdmi_out0_valid_n3 = 1'd0;
reg hdmi_out0_first_n0 = 1'd0;
reg hdmi_out0_last_n0 = 1'd0;
reg hdmi_out0_first_n1 = 1'd0;
reg hdmi_out0_last_n1 = 1'd0;
reg hdmi_out0_first_n2 = 1'd0;
reg hdmi_out0_last_n2 = 1'd0;
reg hdmi_out0_first_n3 = 1'd0;
reg hdmi_out0_last_n3 = 1'd0;
wire hdmi_out0_sink_payload_hsync;
wire hdmi_out0_sink_payload_vsync;
wire hdmi_out0_sink_payload_de;
wire hdmi_out0_source_payload_hsync;
wire hdmi_out0_source_payload_vsync;
wire hdmi_out0_source_payload_de;
reg hdmi_out0_next_s0 = 1'd0;
reg hdmi_out0_next_s1 = 1'd0;
reg hdmi_out0_next_s2 = 1'd0;
reg hdmi_out0_next_s3 = 1'd0;
reg hdmi_out0_next_s4 = 1'd0;
reg hdmi_out0_next_s5 = 1'd0;
reg hdmi_out0_next_s6 = 1'd0;
reg hdmi_out0_next_s7 = 1'd0;
reg hdmi_out0_next_s8 = 1'd0;
reg hdmi_out0_next_s9 = 1'd0;
reg hdmi_out0_next_s10 = 1'd0;
reg hdmi_out0_next_s11 = 1'd0;
reg hdmi_out0_next_s12 = 1'd0;
reg hdmi_out0_next_s13 = 1'd0;
reg hdmi_out0_next_s14 = 1'd0;
reg hdmi_out0_next_s15 = 1'd0;
reg hdmi_out0_next_s16 = 1'd0;
reg hdmi_out0_next_s17 = 1'd0;
reg hdmi_out0_de_r = 1'd0;
reg hdmi_out0_core_source_valid_d = 1'd0;
reg [15:0] hdmi_out0_core_source_data_d = 16'd0;
reg [2:0] wishbonestreamingbridge_state = 3'd0;
reg [2:0] wishbonestreamingbridge_next_state = 3'd0;
reg [1:0] oled_state = 2'd0;
reg [1:0] oled_next_state = 2'd0;
reg [1:0] refresher_state = 2'd0;
reg [1:0] refresher_next_state = 2'd0;
reg [2:0] bankmachine0_state = 3'd0;
reg [2:0] bankmachine0_next_state = 3'd0;
reg [2:0] bankmachine1_state = 3'd0;
reg [2:0] bankmachine1_next_state = 3'd0;
reg [2:0] bankmachine2_state = 3'd0;
reg [2:0] bankmachine2_next_state = 3'd0;
reg [2:0] bankmachine3_state = 3'd0;
reg [2:0] bankmachine3_next_state = 3'd0;
reg [2:0] bankmachine4_state = 3'd0;
reg [2:0] bankmachine4_next_state = 3'd0;
reg [2:0] bankmachine5_state = 3'd0;
reg [2:0] bankmachine5_next_state = 3'd0;
reg [2:0] bankmachine6_state = 3'd0;
reg [2:0] bankmachine6_next_state = 3'd0;
reg [2:0] bankmachine7_state = 3'd0;
reg [2:0] bankmachine7_next_state = 3'd0;
reg [3:0] multiplexer_state = 4'd0;
reg [3:0] multiplexer_next_state = 4'd0;
wire [2:0] cba0;
wire [21:0] rca0;
wire [2:0] cba1;
wire [21:0] rca1;
wire [2:0] cba2;
wire [21:0] rca2;
wire [2:0] roundrobin0_request;
reg [1:0] roundrobin0_grant = 2'd0;
wire roundrobin0_ce;
wire [2:0] roundrobin1_request;
reg [1:0] roundrobin1_grant = 2'd0;
wire roundrobin1_ce;
wire [2:0] roundrobin2_request;
reg [1:0] roundrobin2_grant = 2'd0;
wire roundrobin2_ce;
wire [2:0] roundrobin3_request;
reg [1:0] roundrobin3_grant = 2'd0;
wire roundrobin3_ce;
wire [2:0] roundrobin4_request;
reg [1:0] roundrobin4_grant = 2'd0;
wire roundrobin4_ce;
wire [2:0] roundrobin5_request;
reg [1:0] roundrobin5_grant = 2'd0;
wire roundrobin5_ce;
wire [2:0] roundrobin6_request;
reg [1:0] roundrobin6_grant = 2'd0;
wire roundrobin6_ce;
wire [2:0] roundrobin7_request;
reg [1:0] roundrobin7_grant = 2'd0;
wire roundrobin7_ce;
reg new_master_wdata_ready0 = 1'd0;
reg new_master_wdata_ready1 = 1'd0;
reg new_master_wdata_ready2 = 1'd0;
reg new_master_wdata_ready3 = 1'd0;
reg new_master_wdata_ready4 = 1'd0;
reg new_master_wdata_ready5 = 1'd0;
reg new_master_wdata_ready6 = 1'd0;
reg new_master_wdata_ready7 = 1'd0;
reg new_master_wdata_ready8 = 1'd0;
reg new_master_rdata_valid0 = 1'd0;
reg new_master_rdata_valid1 = 1'd0;
reg new_master_rdata_valid2 = 1'd0;
reg new_master_rdata_valid3 = 1'd0;
reg new_master_rdata_valid4 = 1'd0;
reg new_master_rdata_valid5 = 1'd0;
reg new_master_rdata_valid6 = 1'd0;
reg new_master_rdata_valid7 = 1'd0;
reg new_master_rdata_valid8 = 1'd0;
reg new_master_rdata_valid9 = 1'd0;
reg new_master_rdata_valid10 = 1'd0;
reg new_master_rdata_valid11 = 1'd0;
reg new_master_rdata_valid12 = 1'd0;
reg new_master_rdata_valid13 = 1'd0;
reg new_master_rdata_valid14 = 1'd0;
reg new_master_rdata_valid15 = 1'd0;
reg new_master_rdata_valid16 = 1'd0;
reg new_master_rdata_valid17 = 1'd0;
reg new_master_rdata_valid18 = 1'd0;
reg new_master_rdata_valid19 = 1'd0;
reg new_master_rdata_valid20 = 1'd0;
reg [2:0] fullmemorywe_state = 3'd0;
reg [2:0] fullmemorywe_next_state = 3'd0;
reg [1:0] litedramwishbonebridge_state = 2'd0;
reg [1:0] litedramwishbonebridge_next_state = 2'd0;
reg liteethmacgap_state = 1'd0;
reg liteethmacgap_next_state = 1'd0;
reg [1:0] liteethmacpreambleinserter_state = 2'd0;
reg [1:0] liteethmacpreambleinserter_next_state = 2'd0;
reg liteethmacpreamblechecker_state = 1'd0;
reg liteethmacpreamblechecker_next_state = 1'd0;
reg [1:0] liteethmaccrc32inserter_state = 2'd0;
reg [1:0] liteethmaccrc32inserter_next_state = 2'd0;
reg [1:0] liteethmaccrc32checker_state = 2'd0;
reg [1:0] liteethmaccrc32checker_next_state = 2'd0;
reg liteethmacpaddinginserter_state = 1'd0;
reg liteethmacpaddinginserter_next_state = 1'd0;
reg [2:0] liteethmacsramwriter_state = 3'd0;
reg [2:0] liteethmacsramwriter_next_state = 3'd0;
reg [31:0] ethmac_writer_errors_status_liteethmac_next_value = 32'd0;
reg ethmac_writer_errors_status_liteethmac_next_value_ce = 1'd0;
reg [1:0] liteethmacsramreader_state = 2'd0;
reg [1:0] liteethmacsramreader_next_state = 2'd0;
reg [3:0] edid_state = 4'd0;
reg [3:0] edid_next_state = 4'd0;
reg [1:0] dma_state = 2'd0;
reg [1:0] dma_next_state = 2'd0;
reg videoout_state = 1'd0;
reg videoout_next_state = 1'd0;
reg [27:0] hdmi_out0_core_dmareader_offset_videoout_next_value = 28'd0;
reg hdmi_out0_core_dmareader_offset_videoout_next_value_ce = 1'd0;
wire wb_sdram_con_request;
wire wb_sdram_con_grant;
wire [29:0] videosoc_shared_adr;
wire [31:0] videosoc_shared_dat_w;
wire [31:0] videosoc_shared_dat_r;
wire [3:0] videosoc_shared_sel;
wire videosoc_shared_cyc;
wire videosoc_shared_stb;
wire videosoc_shared_ack;
wire videosoc_shared_we;
wire [2:0] videosoc_shared_cti;
wire [1:0] videosoc_shared_bte;
wire videosoc_shared_err;
wire [2:0] videosoc_request;
reg [1:0] videosoc_grant = 2'd0;
reg [5:0] videosoc_slave_sel = 6'd0;
reg [5:0] videosoc_slave_sel_r = 6'd0;
wire [13:0] videosoc_interface0_bank_bus_adr;
wire videosoc_interface0_bank_bus_we;
wire [7:0] videosoc_interface0_bank_bus_dat_w;
reg [7:0] videosoc_interface0_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank0_dly_sel0_re;
wire [1:0] videosoc_csrbank0_dly_sel0_r;
wire [1:0] videosoc_csrbank0_dly_sel0_w;
wire videosoc_csrbank0_sel;
wire [13:0] videosoc_interface1_bank_bus_adr;
wire videosoc_interface1_bank_bus_we;
wire [7:0] videosoc_interface1_bank_bus_dat_w;
reg [7:0] videosoc_interface1_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank1_sram_writer_slot_re;
wire videosoc_csrbank1_sram_writer_slot_r;
wire videosoc_csrbank1_sram_writer_slot_w;
wire videosoc_csrbank1_sram_writer_length3_re;
wire [7:0] videosoc_csrbank1_sram_writer_length3_r;
wire [7:0] videosoc_csrbank1_sram_writer_length3_w;
wire videosoc_csrbank1_sram_writer_length2_re;
wire [7:0] videosoc_csrbank1_sram_writer_length2_r;
wire [7:0] videosoc_csrbank1_sram_writer_length2_w;
wire videosoc_csrbank1_sram_writer_length1_re;
wire [7:0] videosoc_csrbank1_sram_writer_length1_r;
wire [7:0] videosoc_csrbank1_sram_writer_length1_w;
wire videosoc_csrbank1_sram_writer_length0_re;
wire [7:0] videosoc_csrbank1_sram_writer_length0_r;
wire [7:0] videosoc_csrbank1_sram_writer_length0_w;
wire videosoc_csrbank1_sram_writer_errors3_re;
wire [7:0] videosoc_csrbank1_sram_writer_errors3_r;
wire [7:0] videosoc_csrbank1_sram_writer_errors3_w;
wire videosoc_csrbank1_sram_writer_errors2_re;
wire [7:0] videosoc_csrbank1_sram_writer_errors2_r;
wire [7:0] videosoc_csrbank1_sram_writer_errors2_w;
wire videosoc_csrbank1_sram_writer_errors1_re;
wire [7:0] videosoc_csrbank1_sram_writer_errors1_r;
wire [7:0] videosoc_csrbank1_sram_writer_errors1_w;
wire videosoc_csrbank1_sram_writer_errors0_re;
wire [7:0] videosoc_csrbank1_sram_writer_errors0_r;
wire [7:0] videosoc_csrbank1_sram_writer_errors0_w;
wire videosoc_csrbank1_sram_writer_ev_enable0_re;
wire videosoc_csrbank1_sram_writer_ev_enable0_r;
wire videosoc_csrbank1_sram_writer_ev_enable0_w;
wire videosoc_csrbank1_sram_reader_ready_re;
wire videosoc_csrbank1_sram_reader_ready_r;
wire videosoc_csrbank1_sram_reader_ready_w;
wire videosoc_csrbank1_sram_reader_level_re;
wire [1:0] videosoc_csrbank1_sram_reader_level_r;
wire [1:0] videosoc_csrbank1_sram_reader_level_w;
wire videosoc_csrbank1_sram_reader_slot0_re;
wire videosoc_csrbank1_sram_reader_slot0_r;
wire videosoc_csrbank1_sram_reader_slot0_w;
wire videosoc_csrbank1_sram_reader_length1_re;
wire [2:0] videosoc_csrbank1_sram_reader_length1_r;
wire [2:0] videosoc_csrbank1_sram_reader_length1_w;
wire videosoc_csrbank1_sram_reader_length0_re;
wire [7:0] videosoc_csrbank1_sram_reader_length0_r;
wire [7:0] videosoc_csrbank1_sram_reader_length0_w;
wire videosoc_csrbank1_sram_reader_ev_enable0_re;
wire videosoc_csrbank1_sram_reader_ev_enable0_r;
wire videosoc_csrbank1_sram_reader_ev_enable0_w;
wire videosoc_csrbank1_preamble_crc_re;
wire videosoc_csrbank1_preamble_crc_r;
wire videosoc_csrbank1_preamble_crc_w;
wire videosoc_csrbank1_preamble_errors3_re;
wire [7:0] videosoc_csrbank1_preamble_errors3_r;
wire [7:0] videosoc_csrbank1_preamble_errors3_w;
wire videosoc_csrbank1_preamble_errors2_re;
wire [7:0] videosoc_csrbank1_preamble_errors2_r;
wire [7:0] videosoc_csrbank1_preamble_errors2_w;
wire videosoc_csrbank1_preamble_errors1_re;
wire [7:0] videosoc_csrbank1_preamble_errors1_r;
wire [7:0] videosoc_csrbank1_preamble_errors1_w;
wire videosoc_csrbank1_preamble_errors0_re;
wire [7:0] videosoc_csrbank1_preamble_errors0_r;
wire [7:0] videosoc_csrbank1_preamble_errors0_w;
wire videosoc_csrbank1_crc_errors3_re;
wire [7:0] videosoc_csrbank1_crc_errors3_r;
wire [7:0] videosoc_csrbank1_crc_errors3_w;
wire videosoc_csrbank1_crc_errors2_re;
wire [7:0] videosoc_csrbank1_crc_errors2_r;
wire [7:0] videosoc_csrbank1_crc_errors2_w;
wire videosoc_csrbank1_crc_errors1_re;
wire [7:0] videosoc_csrbank1_crc_errors1_r;
wire [7:0] videosoc_csrbank1_crc_errors1_w;
wire videosoc_csrbank1_crc_errors0_re;
wire [7:0] videosoc_csrbank1_crc_errors0_r;
wire [7:0] videosoc_csrbank1_crc_errors0_w;
wire videosoc_csrbank1_sel;
wire [13:0] videosoc_interface2_bank_bus_adr;
wire videosoc_interface2_bank_bus_we;
wire [7:0] videosoc_interface2_bank_bus_dat_w;
reg [7:0] videosoc_interface2_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank2_crg_reset0_re;
wire videosoc_csrbank2_crg_reset0_r;
wire videosoc_csrbank2_crg_reset0_w;
wire videosoc_csrbank2_mdio_w0_re;
wire [2:0] videosoc_csrbank2_mdio_w0_r;
wire [2:0] videosoc_csrbank2_mdio_w0_w;
wire videosoc_csrbank2_mdio_r_re;
wire videosoc_csrbank2_mdio_r_r;
wire videosoc_csrbank2_mdio_r_w;
wire videosoc_csrbank2_sel;
wire [13:0] videosoc_interface0_sram_bus_adr;
wire videosoc_interface0_sram_bus_we;
wire [7:0] videosoc_interface0_sram_bus_dat_w;
reg [7:0] videosoc_interface0_sram_bus_dat_r = 8'd0;
wire [6:0] videosoc_sram0_adr;
wire [7:0] videosoc_sram0_dat_r;
wire videosoc_sram0_we;
wire [7:0] videosoc_sram0_dat_w;
wire videosoc_sram0_sel;
reg videosoc_sram0_sel_r = 1'd0;
wire [13:0] videosoc_interface3_bank_bus_adr;
wire videosoc_interface3_bank_bus_we;
wire [7:0] videosoc_interface3_bank_bus_dat_w;
reg [7:0] videosoc_interface3_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank3_edid_hpd_notif_re;
wire videosoc_csrbank3_edid_hpd_notif_r;
wire videosoc_csrbank3_edid_hpd_notif_w;
wire videosoc_csrbank3_edid_hpd_en0_re;
wire videosoc_csrbank3_edid_hpd_en0_r;
wire videosoc_csrbank3_edid_hpd_en0_w;
wire videosoc_csrbank3_clocking_mmcm_reset0_re;
wire videosoc_csrbank3_clocking_mmcm_reset0_r;
wire videosoc_csrbank3_clocking_mmcm_reset0_w;
wire videosoc_csrbank3_clocking_locked_re;
wire videosoc_csrbank3_clocking_locked_r;
wire videosoc_csrbank3_clocking_locked_w;
wire videosoc_csrbank3_clocking_mmcm_drdy_re;
wire videosoc_csrbank3_clocking_mmcm_drdy_r;
wire videosoc_csrbank3_clocking_mmcm_drdy_w;
wire videosoc_csrbank3_clocking_mmcm_adr0_re;
wire [6:0] videosoc_csrbank3_clocking_mmcm_adr0_r;
wire [6:0] videosoc_csrbank3_clocking_mmcm_adr0_w;
wire videosoc_csrbank3_clocking_mmcm_dat_w1_re;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_w1_r;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_w1_w;
wire videosoc_csrbank3_clocking_mmcm_dat_w0_re;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_w0_r;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_w0_w;
wire videosoc_csrbank3_clocking_mmcm_dat_r1_re;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_r1_r;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_r1_w;
wire videosoc_csrbank3_clocking_mmcm_dat_r0_re;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_r0_r;
wire [7:0] videosoc_csrbank3_clocking_mmcm_dat_r0_w;
wire videosoc_csrbank3_data0_cap_phase_re;
wire [1:0] videosoc_csrbank3_data0_cap_phase_r;
wire [1:0] videosoc_csrbank3_data0_cap_phase_w;
wire videosoc_csrbank3_data0_charsync_char_synced_re;
wire videosoc_csrbank3_data0_charsync_char_synced_r;
wire videosoc_csrbank3_data0_charsync_char_synced_w;
wire videosoc_csrbank3_data0_charsync_ctl_pos_re;
wire [3:0] videosoc_csrbank3_data0_charsync_ctl_pos_r;
wire [3:0] videosoc_csrbank3_data0_charsync_ctl_pos_w;
wire videosoc_csrbank3_data0_wer_value2_re;
wire [7:0] videosoc_csrbank3_data0_wer_value2_r;
wire [7:0] videosoc_csrbank3_data0_wer_value2_w;
wire videosoc_csrbank3_data0_wer_value1_re;
wire [7:0] videosoc_csrbank3_data0_wer_value1_r;
wire [7:0] videosoc_csrbank3_data0_wer_value1_w;
wire videosoc_csrbank3_data0_wer_value0_re;
wire [7:0] videosoc_csrbank3_data0_wer_value0_r;
wire [7:0] videosoc_csrbank3_data0_wer_value0_w;
wire videosoc_csrbank3_data1_cap_phase_re;
wire [1:0] videosoc_csrbank3_data1_cap_phase_r;
wire [1:0] videosoc_csrbank3_data1_cap_phase_w;
wire videosoc_csrbank3_data1_charsync_char_synced_re;
wire videosoc_csrbank3_data1_charsync_char_synced_r;
wire videosoc_csrbank3_data1_charsync_char_synced_w;
wire videosoc_csrbank3_data1_charsync_ctl_pos_re;
wire [3:0] videosoc_csrbank3_data1_charsync_ctl_pos_r;
wire [3:0] videosoc_csrbank3_data1_charsync_ctl_pos_w;
wire videosoc_csrbank3_data1_wer_value2_re;
wire [7:0] videosoc_csrbank3_data1_wer_value2_r;
wire [7:0] videosoc_csrbank3_data1_wer_value2_w;
wire videosoc_csrbank3_data1_wer_value1_re;
wire [7:0] videosoc_csrbank3_data1_wer_value1_r;
wire [7:0] videosoc_csrbank3_data1_wer_value1_w;
wire videosoc_csrbank3_data1_wer_value0_re;
wire [7:0] videosoc_csrbank3_data1_wer_value0_r;
wire [7:0] videosoc_csrbank3_data1_wer_value0_w;
wire videosoc_csrbank3_data2_cap_phase_re;
wire [1:0] videosoc_csrbank3_data2_cap_phase_r;
wire [1:0] videosoc_csrbank3_data2_cap_phase_w;
wire videosoc_csrbank3_data2_charsync_char_synced_re;
wire videosoc_csrbank3_data2_charsync_char_synced_r;
wire videosoc_csrbank3_data2_charsync_char_synced_w;
wire videosoc_csrbank3_data2_charsync_ctl_pos_re;
wire [3:0] videosoc_csrbank3_data2_charsync_ctl_pos_r;
wire [3:0] videosoc_csrbank3_data2_charsync_ctl_pos_w;
wire videosoc_csrbank3_data2_wer_value2_re;
wire [7:0] videosoc_csrbank3_data2_wer_value2_r;
wire [7:0] videosoc_csrbank3_data2_wer_value2_w;
wire videosoc_csrbank3_data2_wer_value1_re;
wire [7:0] videosoc_csrbank3_data2_wer_value1_r;
wire [7:0] videosoc_csrbank3_data2_wer_value1_w;
wire videosoc_csrbank3_data2_wer_value0_re;
wire [7:0] videosoc_csrbank3_data2_wer_value0_r;
wire [7:0] videosoc_csrbank3_data2_wer_value0_w;
wire videosoc_csrbank3_chansync_channels_synced_re;
wire videosoc_csrbank3_chansync_channels_synced_r;
wire videosoc_csrbank3_chansync_channels_synced_w;
wire videosoc_csrbank3_resdetection_hres1_re;
wire [2:0] videosoc_csrbank3_resdetection_hres1_r;
wire [2:0] videosoc_csrbank3_resdetection_hres1_w;
wire videosoc_csrbank3_resdetection_hres0_re;
wire [7:0] videosoc_csrbank3_resdetection_hres0_r;
wire [7:0] videosoc_csrbank3_resdetection_hres0_w;
wire videosoc_csrbank3_resdetection_vres1_re;
wire [2:0] videosoc_csrbank3_resdetection_vres1_r;
wire [2:0] videosoc_csrbank3_resdetection_vres1_w;
wire videosoc_csrbank3_resdetection_vres0_re;
wire [7:0] videosoc_csrbank3_resdetection_vres0_r;
wire [7:0] videosoc_csrbank3_resdetection_vres0_w;
wire videosoc_csrbank3_dma_frame_size3_re;
wire [4:0] videosoc_csrbank3_dma_frame_size3_r;
wire [4:0] videosoc_csrbank3_dma_frame_size3_w;
wire videosoc_csrbank3_dma_frame_size2_re;
wire [7:0] videosoc_csrbank3_dma_frame_size2_r;
wire [7:0] videosoc_csrbank3_dma_frame_size2_w;
wire videosoc_csrbank3_dma_frame_size1_re;
wire [7:0] videosoc_csrbank3_dma_frame_size1_r;
wire [7:0] videosoc_csrbank3_dma_frame_size1_w;
wire videosoc_csrbank3_dma_frame_size0_re;
wire [7:0] videosoc_csrbank3_dma_frame_size0_r;
wire [7:0] videosoc_csrbank3_dma_frame_size0_w;
wire videosoc_csrbank3_dma_slot0_status0_re;
wire [1:0] videosoc_csrbank3_dma_slot0_status0_r;
wire [1:0] videosoc_csrbank3_dma_slot0_status0_w;
wire videosoc_csrbank3_dma_slot0_address3_re;
wire [4:0] videosoc_csrbank3_dma_slot0_address3_r;
wire [4:0] videosoc_csrbank3_dma_slot0_address3_w;
wire videosoc_csrbank3_dma_slot0_address2_re;
wire [7:0] videosoc_csrbank3_dma_slot0_address2_r;
wire [7:0] videosoc_csrbank3_dma_slot0_address2_w;
wire videosoc_csrbank3_dma_slot0_address1_re;
wire [7:0] videosoc_csrbank3_dma_slot0_address1_r;
wire [7:0] videosoc_csrbank3_dma_slot0_address1_w;
wire videosoc_csrbank3_dma_slot0_address0_re;
wire [7:0] videosoc_csrbank3_dma_slot0_address0_r;
wire [7:0] videosoc_csrbank3_dma_slot0_address0_w;
wire videosoc_csrbank3_dma_slot1_status0_re;
wire [1:0] videosoc_csrbank3_dma_slot1_status0_r;
wire [1:0] videosoc_csrbank3_dma_slot1_status0_w;
wire videosoc_csrbank3_dma_slot1_address3_re;
wire [4:0] videosoc_csrbank3_dma_slot1_address3_r;
wire [4:0] videosoc_csrbank3_dma_slot1_address3_w;
wire videosoc_csrbank3_dma_slot1_address2_re;
wire [7:0] videosoc_csrbank3_dma_slot1_address2_r;
wire [7:0] videosoc_csrbank3_dma_slot1_address2_w;
wire videosoc_csrbank3_dma_slot1_address1_re;
wire [7:0] videosoc_csrbank3_dma_slot1_address1_r;
wire [7:0] videosoc_csrbank3_dma_slot1_address1_w;
wire videosoc_csrbank3_dma_slot1_address0_re;
wire [7:0] videosoc_csrbank3_dma_slot1_address0_r;
wire [7:0] videosoc_csrbank3_dma_slot1_address0_w;
wire videosoc_csrbank3_dma_ev_enable0_re;
wire [1:0] videosoc_csrbank3_dma_ev_enable0_r;
wire [1:0] videosoc_csrbank3_dma_ev_enable0_w;
wire videosoc_csrbank3_sel;
wire [13:0] videosoc_interface4_bank_bus_adr;
wire videosoc_interface4_bank_bus_we;
wire [7:0] videosoc_interface4_bank_bus_dat_w;
reg [7:0] videosoc_interface4_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank4_value3_re;
wire [7:0] videosoc_csrbank4_value3_r;
wire [7:0] videosoc_csrbank4_value3_w;
wire videosoc_csrbank4_value2_re;
wire [7:0] videosoc_csrbank4_value2_r;
wire [7:0] videosoc_csrbank4_value2_w;
wire videosoc_csrbank4_value1_re;
wire [7:0] videosoc_csrbank4_value1_r;
wire [7:0] videosoc_csrbank4_value1_w;
wire videosoc_csrbank4_value0_re;
wire [7:0] videosoc_csrbank4_value0_r;
wire [7:0] videosoc_csrbank4_value0_w;
wire videosoc_csrbank4_sel;
wire [13:0] videosoc_interface5_bank_bus_adr;
wire videosoc_interface5_bank_bus_we;
wire [7:0] videosoc_interface5_bank_bus_dat_w;
reg [7:0] videosoc_interface5_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank5_core_underflow_enable0_re;
wire videosoc_csrbank5_core_underflow_enable0_r;
wire videosoc_csrbank5_core_underflow_enable0_w;
wire videosoc_csrbank5_core_underflow_counter3_re;
wire [7:0] videosoc_csrbank5_core_underflow_counter3_r;
wire [7:0] videosoc_csrbank5_core_underflow_counter3_w;
wire videosoc_csrbank5_core_underflow_counter2_re;
wire [7:0] videosoc_csrbank5_core_underflow_counter2_r;
wire [7:0] videosoc_csrbank5_core_underflow_counter2_w;
wire videosoc_csrbank5_core_underflow_counter1_re;
wire [7:0] videosoc_csrbank5_core_underflow_counter1_r;
wire [7:0] videosoc_csrbank5_core_underflow_counter1_w;
wire videosoc_csrbank5_core_underflow_counter0_re;
wire [7:0] videosoc_csrbank5_core_underflow_counter0_r;
wire [7:0] videosoc_csrbank5_core_underflow_counter0_w;
wire videosoc_csrbank5_core_initiator_enable0_re;
wire videosoc_csrbank5_core_initiator_enable0_r;
wire videosoc_csrbank5_core_initiator_enable0_w;
reg [3:0] videosoc_csrbank5_core_initiator_hres_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_hres1_re;
wire [3:0] videosoc_csrbank5_core_initiator_hres1_r;
wire [3:0] videosoc_csrbank5_core_initiator_hres1_w;
wire videosoc_csrbank5_core_initiator_hres0_re;
wire [7:0] videosoc_csrbank5_core_initiator_hres0_r;
wire [7:0] videosoc_csrbank5_core_initiator_hres0_w;
reg [3:0] videosoc_csrbank5_core_initiator_hsync_start_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_hsync_start1_re;
wire [3:0] videosoc_csrbank5_core_initiator_hsync_start1_r;
wire [3:0] videosoc_csrbank5_core_initiator_hsync_start1_w;
wire videosoc_csrbank5_core_initiator_hsync_start0_re;
wire [7:0] videosoc_csrbank5_core_initiator_hsync_start0_r;
wire [7:0] videosoc_csrbank5_core_initiator_hsync_start0_w;
reg [3:0] videosoc_csrbank5_core_initiator_hsync_end_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_hsync_end1_re;
wire [3:0] videosoc_csrbank5_core_initiator_hsync_end1_r;
wire [3:0] videosoc_csrbank5_core_initiator_hsync_end1_w;
wire videosoc_csrbank5_core_initiator_hsync_end0_re;
wire [7:0] videosoc_csrbank5_core_initiator_hsync_end0_r;
wire [7:0] videosoc_csrbank5_core_initiator_hsync_end0_w;
reg [3:0] videosoc_csrbank5_core_initiator_hscan_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_hscan1_re;
wire [3:0] videosoc_csrbank5_core_initiator_hscan1_r;
wire [3:0] videosoc_csrbank5_core_initiator_hscan1_w;
wire videosoc_csrbank5_core_initiator_hscan0_re;
wire [7:0] videosoc_csrbank5_core_initiator_hscan0_r;
wire [7:0] videosoc_csrbank5_core_initiator_hscan0_w;
reg [3:0] videosoc_csrbank5_core_initiator_vres_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_vres1_re;
wire [3:0] videosoc_csrbank5_core_initiator_vres1_r;
wire [3:0] videosoc_csrbank5_core_initiator_vres1_w;
wire videosoc_csrbank5_core_initiator_vres0_re;
wire [7:0] videosoc_csrbank5_core_initiator_vres0_r;
wire [7:0] videosoc_csrbank5_core_initiator_vres0_w;
reg [3:0] videosoc_csrbank5_core_initiator_vsync_start_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_vsync_start1_re;
wire [3:0] videosoc_csrbank5_core_initiator_vsync_start1_r;
wire [3:0] videosoc_csrbank5_core_initiator_vsync_start1_w;
wire videosoc_csrbank5_core_initiator_vsync_start0_re;
wire [7:0] videosoc_csrbank5_core_initiator_vsync_start0_r;
wire [7:0] videosoc_csrbank5_core_initiator_vsync_start0_w;
reg [3:0] videosoc_csrbank5_core_initiator_vsync_end_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_vsync_end1_re;
wire [3:0] videosoc_csrbank5_core_initiator_vsync_end1_r;
wire [3:0] videosoc_csrbank5_core_initiator_vsync_end1_w;
wire videosoc_csrbank5_core_initiator_vsync_end0_re;
wire [7:0] videosoc_csrbank5_core_initiator_vsync_end0_r;
wire [7:0] videosoc_csrbank5_core_initiator_vsync_end0_w;
reg [3:0] videosoc_csrbank5_core_initiator_vscan_backstore = 4'd0;
wire videosoc_csrbank5_core_initiator_vscan1_re;
wire [3:0] videosoc_csrbank5_core_initiator_vscan1_r;
wire [3:0] videosoc_csrbank5_core_initiator_vscan1_w;
wire videosoc_csrbank5_core_initiator_vscan0_re;
wire [7:0] videosoc_csrbank5_core_initiator_vscan0_r;
wire [7:0] videosoc_csrbank5_core_initiator_vscan0_w;
reg [23:0] videosoc_csrbank5_core_initiator_base_backstore = 24'd0;
wire videosoc_csrbank5_core_initiator_base3_re;
wire [7:0] videosoc_csrbank5_core_initiator_base3_r;
wire [7:0] videosoc_csrbank5_core_initiator_base3_w;
wire videosoc_csrbank5_core_initiator_base2_re;
wire [7:0] videosoc_csrbank5_core_initiator_base2_r;
wire [7:0] videosoc_csrbank5_core_initiator_base2_w;
wire videosoc_csrbank5_core_initiator_base1_re;
wire [7:0] videosoc_csrbank5_core_initiator_base1_r;
wire [7:0] videosoc_csrbank5_core_initiator_base1_w;
wire videosoc_csrbank5_core_initiator_base0_re;
wire [7:0] videosoc_csrbank5_core_initiator_base0_r;
wire [7:0] videosoc_csrbank5_core_initiator_base0_w;
reg [23:0] videosoc_csrbank5_core_initiator_length_backstore = 24'd0;
wire videosoc_csrbank5_core_initiator_length3_re;
wire [7:0] videosoc_csrbank5_core_initiator_length3_r;
wire [7:0] videosoc_csrbank5_core_initiator_length3_w;
wire videosoc_csrbank5_core_initiator_length2_re;
wire [7:0] videosoc_csrbank5_core_initiator_length2_r;
wire [7:0] videosoc_csrbank5_core_initiator_length2_w;
wire videosoc_csrbank5_core_initiator_length1_re;
wire [7:0] videosoc_csrbank5_core_initiator_length1_r;
wire [7:0] videosoc_csrbank5_core_initiator_length1_w;
wire videosoc_csrbank5_core_initiator_length0_re;
wire [7:0] videosoc_csrbank5_core_initiator_length0_r;
wire [7:0] videosoc_csrbank5_core_initiator_length0_w;
wire videosoc_csrbank5_driver_clocking_mmcm_reset0_re;
wire videosoc_csrbank5_driver_clocking_mmcm_reset0_r;
wire videosoc_csrbank5_driver_clocking_mmcm_reset0_w;
wire videosoc_csrbank5_driver_clocking_mmcm_drdy_re;
wire videosoc_csrbank5_driver_clocking_mmcm_drdy_r;
wire videosoc_csrbank5_driver_clocking_mmcm_drdy_w;
wire videosoc_csrbank5_driver_clocking_mmcm_adr0_re;
wire [6:0] videosoc_csrbank5_driver_clocking_mmcm_adr0_r;
wire [6:0] videosoc_csrbank5_driver_clocking_mmcm_adr0_w;
wire videosoc_csrbank5_driver_clocking_mmcm_dat_w1_re;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_w1_r;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_w1_w;
wire videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_w0_r;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_w0_w;
wire videosoc_csrbank5_driver_clocking_mmcm_dat_r1_re;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_r1_r;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_r1_w;
wire videosoc_csrbank5_driver_clocking_mmcm_dat_r0_re;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_r0_r;
wire [7:0] videosoc_csrbank5_driver_clocking_mmcm_dat_r0_w;
wire videosoc_csrbank5_sel;
wire [13:0] videosoc_interface1_sram_bus_adr;
wire videosoc_interface1_sram_bus_we;
wire [7:0] videosoc_interface1_sram_bus_dat_w;
reg [7:0] videosoc_interface1_sram_bus_dat_r = 8'd0;
wire [3:0] videosoc_sram1_adr;
wire [7:0] videosoc_sram1_dat_r;
wire videosoc_sram1_sel;
reg videosoc_sram1_sel_r = 1'd0;
wire [13:0] videosoc_interface6_bank_bus_adr;
wire videosoc_interface6_bank_bus_we;
wire [7:0] videosoc_interface6_bank_bus_dat_w;
reg [7:0] videosoc_interface6_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank6_dna_id7_re;
wire videosoc_csrbank6_dna_id7_r;
wire videosoc_csrbank6_dna_id7_w;
wire videosoc_csrbank6_dna_id6_re;
wire [7:0] videosoc_csrbank6_dna_id6_r;
wire [7:0] videosoc_csrbank6_dna_id6_w;
wire videosoc_csrbank6_dna_id5_re;
wire [7:0] videosoc_csrbank6_dna_id5_r;
wire [7:0] videosoc_csrbank6_dna_id5_w;
wire videosoc_csrbank6_dna_id4_re;
wire [7:0] videosoc_csrbank6_dna_id4_r;
wire [7:0] videosoc_csrbank6_dna_id4_w;
wire videosoc_csrbank6_dna_id3_re;
wire [7:0] videosoc_csrbank6_dna_id3_r;
wire [7:0] videosoc_csrbank6_dna_id3_w;
wire videosoc_csrbank6_dna_id2_re;
wire [7:0] videosoc_csrbank6_dna_id2_r;
wire [7:0] videosoc_csrbank6_dna_id2_w;
wire videosoc_csrbank6_dna_id1_re;
wire [7:0] videosoc_csrbank6_dna_id1_r;
wire [7:0] videosoc_csrbank6_dna_id1_w;
wire videosoc_csrbank6_dna_id0_re;
wire [7:0] videosoc_csrbank6_dna_id0_r;
wire [7:0] videosoc_csrbank6_dna_id0_w;
wire videosoc_csrbank6_git_commit19_re;
wire [7:0] videosoc_csrbank6_git_commit19_r;
wire [7:0] videosoc_csrbank6_git_commit19_w;
wire videosoc_csrbank6_git_commit18_re;
wire [7:0] videosoc_csrbank6_git_commit18_r;
wire [7:0] videosoc_csrbank6_git_commit18_w;
wire videosoc_csrbank6_git_commit17_re;
wire [7:0] videosoc_csrbank6_git_commit17_r;
wire [7:0] videosoc_csrbank6_git_commit17_w;
wire videosoc_csrbank6_git_commit16_re;
wire [7:0] videosoc_csrbank6_git_commit16_r;
wire [7:0] videosoc_csrbank6_git_commit16_w;
wire videosoc_csrbank6_git_commit15_re;
wire [7:0] videosoc_csrbank6_git_commit15_r;
wire [7:0] videosoc_csrbank6_git_commit15_w;
wire videosoc_csrbank6_git_commit14_re;
wire [7:0] videosoc_csrbank6_git_commit14_r;
wire [7:0] videosoc_csrbank6_git_commit14_w;
wire videosoc_csrbank6_git_commit13_re;
wire [7:0] videosoc_csrbank6_git_commit13_r;
wire [7:0] videosoc_csrbank6_git_commit13_w;
wire videosoc_csrbank6_git_commit12_re;
wire [7:0] videosoc_csrbank6_git_commit12_r;
wire [7:0] videosoc_csrbank6_git_commit12_w;
wire videosoc_csrbank6_git_commit11_re;
wire [7:0] videosoc_csrbank6_git_commit11_r;
wire [7:0] videosoc_csrbank6_git_commit11_w;
wire videosoc_csrbank6_git_commit10_re;
wire [7:0] videosoc_csrbank6_git_commit10_r;
wire [7:0] videosoc_csrbank6_git_commit10_w;
wire videosoc_csrbank6_git_commit9_re;
wire [7:0] videosoc_csrbank6_git_commit9_r;
wire [7:0] videosoc_csrbank6_git_commit9_w;
wire videosoc_csrbank6_git_commit8_re;
wire [7:0] videosoc_csrbank6_git_commit8_r;
wire [7:0] videosoc_csrbank6_git_commit8_w;
wire videosoc_csrbank6_git_commit7_re;
wire [7:0] videosoc_csrbank6_git_commit7_r;
wire [7:0] videosoc_csrbank6_git_commit7_w;
wire videosoc_csrbank6_git_commit6_re;
wire [7:0] videosoc_csrbank6_git_commit6_r;
wire [7:0] videosoc_csrbank6_git_commit6_w;
wire videosoc_csrbank6_git_commit5_re;
wire [7:0] videosoc_csrbank6_git_commit5_r;
wire [7:0] videosoc_csrbank6_git_commit5_w;
wire videosoc_csrbank6_git_commit4_re;
wire [7:0] videosoc_csrbank6_git_commit4_r;
wire [7:0] videosoc_csrbank6_git_commit4_w;
wire videosoc_csrbank6_git_commit3_re;
wire [7:0] videosoc_csrbank6_git_commit3_r;
wire [7:0] videosoc_csrbank6_git_commit3_w;
wire videosoc_csrbank6_git_commit2_re;
wire [7:0] videosoc_csrbank6_git_commit2_r;
wire [7:0] videosoc_csrbank6_git_commit2_w;
wire videosoc_csrbank6_git_commit1_re;
wire [7:0] videosoc_csrbank6_git_commit1_r;
wire [7:0] videosoc_csrbank6_git_commit1_w;
wire videosoc_csrbank6_git_commit0_re;
wire [7:0] videosoc_csrbank6_git_commit0_r;
wire [7:0] videosoc_csrbank6_git_commit0_w;
wire videosoc_csrbank6_platform_platform7_re;
wire [7:0] videosoc_csrbank6_platform_platform7_r;
wire [7:0] videosoc_csrbank6_platform_platform7_w;
wire videosoc_csrbank6_platform_platform6_re;
wire [7:0] videosoc_csrbank6_platform_platform6_r;
wire [7:0] videosoc_csrbank6_platform_platform6_w;
wire videosoc_csrbank6_platform_platform5_re;
wire [7:0] videosoc_csrbank6_platform_platform5_r;
wire [7:0] videosoc_csrbank6_platform_platform5_w;
wire videosoc_csrbank6_platform_platform4_re;
wire [7:0] videosoc_csrbank6_platform_platform4_r;
wire [7:0] videosoc_csrbank6_platform_platform4_w;
wire videosoc_csrbank6_platform_platform3_re;
wire [7:0] videosoc_csrbank6_platform_platform3_r;
wire [7:0] videosoc_csrbank6_platform_platform3_w;
wire videosoc_csrbank6_platform_platform2_re;
wire [7:0] videosoc_csrbank6_platform_platform2_r;
wire [7:0] videosoc_csrbank6_platform_platform2_w;
wire videosoc_csrbank6_platform_platform1_re;
wire [7:0] videosoc_csrbank6_platform_platform1_r;
wire [7:0] videosoc_csrbank6_platform_platform1_w;
wire videosoc_csrbank6_platform_platform0_re;
wire [7:0] videosoc_csrbank6_platform_platform0_r;
wire [7:0] videosoc_csrbank6_platform_platform0_w;
wire videosoc_csrbank6_platform_target7_re;
wire [7:0] videosoc_csrbank6_platform_target7_r;
wire [7:0] videosoc_csrbank6_platform_target7_w;
wire videosoc_csrbank6_platform_target6_re;
wire [7:0] videosoc_csrbank6_platform_target6_r;
wire [7:0] videosoc_csrbank6_platform_target6_w;
wire videosoc_csrbank6_platform_target5_re;
wire [7:0] videosoc_csrbank6_platform_target5_r;
wire [7:0] videosoc_csrbank6_platform_target5_w;
wire videosoc_csrbank6_platform_target4_re;
wire [7:0] videosoc_csrbank6_platform_target4_r;
wire [7:0] videosoc_csrbank6_platform_target4_w;
wire videosoc_csrbank6_platform_target3_re;
wire [7:0] videosoc_csrbank6_platform_target3_r;
wire [7:0] videosoc_csrbank6_platform_target3_w;
wire videosoc_csrbank6_platform_target2_re;
wire [7:0] videosoc_csrbank6_platform_target2_r;
wire [7:0] videosoc_csrbank6_platform_target2_w;
wire videosoc_csrbank6_platform_target1_re;
wire [7:0] videosoc_csrbank6_platform_target1_r;
wire [7:0] videosoc_csrbank6_platform_target1_w;
wire videosoc_csrbank6_platform_target0_re;
wire [7:0] videosoc_csrbank6_platform_target0_r;
wire [7:0] videosoc_csrbank6_platform_target0_w;
wire videosoc_csrbank6_xadc_temperature1_re;
wire [3:0] videosoc_csrbank6_xadc_temperature1_r;
wire [3:0] videosoc_csrbank6_xadc_temperature1_w;
wire videosoc_csrbank6_xadc_temperature0_re;
wire [7:0] videosoc_csrbank6_xadc_temperature0_r;
wire [7:0] videosoc_csrbank6_xadc_temperature0_w;
wire videosoc_csrbank6_xadc_vccint1_re;
wire [3:0] videosoc_csrbank6_xadc_vccint1_r;
wire [3:0] videosoc_csrbank6_xadc_vccint1_w;
wire videosoc_csrbank6_xadc_vccint0_re;
wire [7:0] videosoc_csrbank6_xadc_vccint0_r;
wire [7:0] videosoc_csrbank6_xadc_vccint0_w;
wire videosoc_csrbank6_xadc_vccaux1_re;
wire [3:0] videosoc_csrbank6_xadc_vccaux1_r;
wire [3:0] videosoc_csrbank6_xadc_vccaux1_w;
wire videosoc_csrbank6_xadc_vccaux0_re;
wire [7:0] videosoc_csrbank6_xadc_vccaux0_r;
wire [7:0] videosoc_csrbank6_xadc_vccaux0_w;
wire videosoc_csrbank6_xadc_vccbram1_re;
wire [3:0] videosoc_csrbank6_xadc_vccbram1_r;
wire [3:0] videosoc_csrbank6_xadc_vccbram1_w;
wire videosoc_csrbank6_xadc_vccbram0_re;
wire [7:0] videosoc_csrbank6_xadc_vccbram0_r;
wire [7:0] videosoc_csrbank6_xadc_vccbram0_w;
wire videosoc_csrbank6_sel;
wire [13:0] videosoc_interface7_bank_bus_adr;
wire videosoc_interface7_bank_bus_we;
wire [7:0] videosoc_interface7_bank_bus_dat_w;
reg [7:0] videosoc_interface7_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank7_spi_length0_re;
wire [7:0] videosoc_csrbank7_spi_length0_r;
wire [7:0] videosoc_csrbank7_spi_length0_w;
wire videosoc_csrbank7_spi_status_re;
wire videosoc_csrbank7_spi_status_r;
wire videosoc_csrbank7_spi_status_w;
wire videosoc_csrbank7_spi_mosi0_re;
wire [7:0] videosoc_csrbank7_spi_mosi0_r;
wire [7:0] videosoc_csrbank7_spi_mosi0_w;
wire videosoc_csrbank7_gpio_out0_re;
wire [3:0] videosoc_csrbank7_gpio_out0_r;
wire [3:0] videosoc_csrbank7_gpio_out0_w;
wire videosoc_csrbank7_sel;
wire [13:0] videosoc_interface8_bank_bus_adr;
wire videosoc_interface8_bank_bus_we;
wire [7:0] videosoc_interface8_bank_bus_dat_w;
reg [7:0] videosoc_interface8_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank8_dfii_control0_re;
wire [3:0] videosoc_csrbank8_dfii_control0_r;
wire [3:0] videosoc_csrbank8_dfii_control0_w;
wire videosoc_csrbank8_dfii_pi0_command0_re;
wire [5:0] videosoc_csrbank8_dfii_pi0_command0_r;
wire [5:0] videosoc_csrbank8_dfii_pi0_command0_w;
wire videosoc_csrbank8_dfii_pi0_address1_re;
wire [6:0] videosoc_csrbank8_dfii_pi0_address1_r;
wire [6:0] videosoc_csrbank8_dfii_pi0_address1_w;
wire videosoc_csrbank8_dfii_pi0_address0_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_address0_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_address0_w;
wire videosoc_csrbank8_dfii_pi0_baddress0_re;
wire [2:0] videosoc_csrbank8_dfii_pi0_baddress0_r;
wire [2:0] videosoc_csrbank8_dfii_pi0_baddress0_w;
wire videosoc_csrbank8_dfii_pi0_wrdata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata3_w;
wire videosoc_csrbank8_dfii_pi0_wrdata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata2_w;
wire videosoc_csrbank8_dfii_pi0_wrdata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata1_w;
wire videosoc_csrbank8_dfii_pi0_wrdata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_wrdata0_w;
wire videosoc_csrbank8_dfii_pi0_rddata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata3_w;
wire videosoc_csrbank8_dfii_pi0_rddata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata2_w;
wire videosoc_csrbank8_dfii_pi0_rddata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata1_w;
wire videosoc_csrbank8_dfii_pi0_rddata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi0_rddata0_w;
wire videosoc_csrbank8_dfii_pi1_command0_re;
wire [5:0] videosoc_csrbank8_dfii_pi1_command0_r;
wire [5:0] videosoc_csrbank8_dfii_pi1_command0_w;
wire videosoc_csrbank8_dfii_pi1_address1_re;
wire [6:0] videosoc_csrbank8_dfii_pi1_address1_r;
wire [6:0] videosoc_csrbank8_dfii_pi1_address1_w;
wire videosoc_csrbank8_dfii_pi1_address0_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_address0_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_address0_w;
wire videosoc_csrbank8_dfii_pi1_baddress0_re;
wire [2:0] videosoc_csrbank8_dfii_pi1_baddress0_r;
wire [2:0] videosoc_csrbank8_dfii_pi1_baddress0_w;
wire videosoc_csrbank8_dfii_pi1_wrdata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata3_w;
wire videosoc_csrbank8_dfii_pi1_wrdata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata2_w;
wire videosoc_csrbank8_dfii_pi1_wrdata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata1_w;
wire videosoc_csrbank8_dfii_pi1_wrdata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_wrdata0_w;
wire videosoc_csrbank8_dfii_pi1_rddata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata3_w;
wire videosoc_csrbank8_dfii_pi1_rddata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata2_w;
wire videosoc_csrbank8_dfii_pi1_rddata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata1_w;
wire videosoc_csrbank8_dfii_pi1_rddata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi1_rddata0_w;
wire videosoc_csrbank8_dfii_pi2_command0_re;
wire [5:0] videosoc_csrbank8_dfii_pi2_command0_r;
wire [5:0] videosoc_csrbank8_dfii_pi2_command0_w;
wire videosoc_csrbank8_dfii_pi2_address1_re;
wire [6:0] videosoc_csrbank8_dfii_pi2_address1_r;
wire [6:0] videosoc_csrbank8_dfii_pi2_address1_w;
wire videosoc_csrbank8_dfii_pi2_address0_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_address0_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_address0_w;
wire videosoc_csrbank8_dfii_pi2_baddress0_re;
wire [2:0] videosoc_csrbank8_dfii_pi2_baddress0_r;
wire [2:0] videosoc_csrbank8_dfii_pi2_baddress0_w;
wire videosoc_csrbank8_dfii_pi2_wrdata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata3_w;
wire videosoc_csrbank8_dfii_pi2_wrdata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata2_w;
wire videosoc_csrbank8_dfii_pi2_wrdata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata1_w;
wire videosoc_csrbank8_dfii_pi2_wrdata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_wrdata0_w;
wire videosoc_csrbank8_dfii_pi2_rddata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata3_w;
wire videosoc_csrbank8_dfii_pi2_rddata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata2_w;
wire videosoc_csrbank8_dfii_pi2_rddata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata1_w;
wire videosoc_csrbank8_dfii_pi2_rddata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi2_rddata0_w;
wire videosoc_csrbank8_dfii_pi3_command0_re;
wire [5:0] videosoc_csrbank8_dfii_pi3_command0_r;
wire [5:0] videosoc_csrbank8_dfii_pi3_command0_w;
wire videosoc_csrbank8_dfii_pi3_address1_re;
wire [6:0] videosoc_csrbank8_dfii_pi3_address1_r;
wire [6:0] videosoc_csrbank8_dfii_pi3_address1_w;
wire videosoc_csrbank8_dfii_pi3_address0_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_address0_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_address0_w;
wire videosoc_csrbank8_dfii_pi3_baddress0_re;
wire [2:0] videosoc_csrbank8_dfii_pi3_baddress0_r;
wire [2:0] videosoc_csrbank8_dfii_pi3_baddress0_w;
wire videosoc_csrbank8_dfii_pi3_wrdata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata3_w;
wire videosoc_csrbank8_dfii_pi3_wrdata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata2_w;
wire videosoc_csrbank8_dfii_pi3_wrdata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata1_w;
wire videosoc_csrbank8_dfii_pi3_wrdata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_wrdata0_w;
wire videosoc_csrbank8_dfii_pi3_rddata3_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata3_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata3_w;
wire videosoc_csrbank8_dfii_pi3_rddata2_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata2_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata2_w;
wire videosoc_csrbank8_dfii_pi3_rddata1_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata1_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata1_w;
wire videosoc_csrbank8_dfii_pi3_rddata0_re;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata0_r;
wire [7:0] videosoc_csrbank8_dfii_pi3_rddata0_w;
wire videosoc_csrbank8_controller_bandwidth_nreads2_re;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nreads2_r;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nreads2_w;
wire videosoc_csrbank8_controller_bandwidth_nreads1_re;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nreads1_r;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nreads1_w;
wire videosoc_csrbank8_controller_bandwidth_nreads0_re;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nreads0_r;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nreads0_w;
wire videosoc_csrbank8_controller_bandwidth_nwrites2_re;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nwrites2_r;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nwrites2_w;
wire videosoc_csrbank8_controller_bandwidth_nwrites1_re;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nwrites1_r;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nwrites1_w;
wire videosoc_csrbank8_controller_bandwidth_nwrites0_re;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nwrites0_r;
wire [7:0] videosoc_csrbank8_controller_bandwidth_nwrites0_w;
wire videosoc_csrbank8_controller_bandwidth_data_width_re;
wire [7:0] videosoc_csrbank8_controller_bandwidth_data_width_r;
wire [7:0] videosoc_csrbank8_controller_bandwidth_data_width_w;
wire videosoc_csrbank8_sel;
wire [13:0] videosoc_interface9_bank_bus_adr;
wire videosoc_interface9_bank_bus_we;
wire [7:0] videosoc_interface9_bank_bus_dat_w;
reg [7:0] videosoc_interface9_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank9_bitbang0_re;
wire [3:0] videosoc_csrbank9_bitbang0_r;
wire [3:0] videosoc_csrbank9_bitbang0_w;
wire videosoc_csrbank9_miso_re;
wire videosoc_csrbank9_miso_r;
wire videosoc_csrbank9_miso_w;
wire videosoc_csrbank9_bitbang_en0_re;
wire videosoc_csrbank9_bitbang_en0_r;
wire videosoc_csrbank9_bitbang_en0_w;
wire videosoc_csrbank9_sel;
wire [13:0] videosoc_interface10_bank_bus_adr;
wire videosoc_interface10_bank_bus_we;
wire [7:0] videosoc_interface10_bank_bus_dat_w;
reg [7:0] videosoc_interface10_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank10_load3_re;
wire [7:0] videosoc_csrbank10_load3_r;
wire [7:0] videosoc_csrbank10_load3_w;
wire videosoc_csrbank10_load2_re;
wire [7:0] videosoc_csrbank10_load2_r;
wire [7:0] videosoc_csrbank10_load2_w;
wire videosoc_csrbank10_load1_re;
wire [7:0] videosoc_csrbank10_load1_r;
wire [7:0] videosoc_csrbank10_load1_w;
wire videosoc_csrbank10_load0_re;
wire [7:0] videosoc_csrbank10_load0_r;
wire [7:0] videosoc_csrbank10_load0_w;
wire videosoc_csrbank10_reload3_re;
wire [7:0] videosoc_csrbank10_reload3_r;
wire [7:0] videosoc_csrbank10_reload3_w;
wire videosoc_csrbank10_reload2_re;
wire [7:0] videosoc_csrbank10_reload2_r;
wire [7:0] videosoc_csrbank10_reload2_w;
wire videosoc_csrbank10_reload1_re;
wire [7:0] videosoc_csrbank10_reload1_r;
wire [7:0] videosoc_csrbank10_reload1_w;
wire videosoc_csrbank10_reload0_re;
wire [7:0] videosoc_csrbank10_reload0_r;
wire [7:0] videosoc_csrbank10_reload0_w;
wire videosoc_csrbank10_en0_re;
wire videosoc_csrbank10_en0_r;
wire videosoc_csrbank10_en0_w;
wire videosoc_csrbank10_value3_re;
wire [7:0] videosoc_csrbank10_value3_r;
wire [7:0] videosoc_csrbank10_value3_w;
wire videosoc_csrbank10_value2_re;
wire [7:0] videosoc_csrbank10_value2_r;
wire [7:0] videosoc_csrbank10_value2_w;
wire videosoc_csrbank10_value1_re;
wire [7:0] videosoc_csrbank10_value1_r;
wire [7:0] videosoc_csrbank10_value1_w;
wire videosoc_csrbank10_value0_re;
wire [7:0] videosoc_csrbank10_value0_r;
wire [7:0] videosoc_csrbank10_value0_w;
wire videosoc_csrbank10_ev_enable0_re;
wire videosoc_csrbank10_ev_enable0_r;
wire videosoc_csrbank10_ev_enable0_w;
wire videosoc_csrbank10_sel;
wire [13:0] videosoc_interface11_bank_bus_adr;
wire videosoc_interface11_bank_bus_we;
wire [7:0] videosoc_interface11_bank_bus_dat_w;
reg [7:0] videosoc_interface11_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank11_txfull_re;
wire videosoc_csrbank11_txfull_r;
wire videosoc_csrbank11_txfull_w;
wire videosoc_csrbank11_rxempty_re;
wire videosoc_csrbank11_rxempty_r;
wire videosoc_csrbank11_rxempty_w;
wire videosoc_csrbank11_ev_enable0_re;
wire [1:0] videosoc_csrbank11_ev_enable0_r;
wire [1:0] videosoc_csrbank11_ev_enable0_w;
wire videosoc_csrbank11_sel;
wire [13:0] videosoc_interface12_bank_bus_adr;
wire videosoc_interface12_bank_bus_we;
wire [7:0] videosoc_interface12_bank_bus_dat_w;
reg [7:0] videosoc_interface12_bank_bus_dat_r = 8'd0;
wire videosoc_csrbank12_tuning_word3_re;
wire [7:0] videosoc_csrbank12_tuning_word3_r;
wire [7:0] videosoc_csrbank12_tuning_word3_w;
wire videosoc_csrbank12_tuning_word2_re;
wire [7:0] videosoc_csrbank12_tuning_word2_r;
wire [7:0] videosoc_csrbank12_tuning_word2_w;
wire videosoc_csrbank12_tuning_word1_re;
wire [7:0] videosoc_csrbank12_tuning_word1_r;
wire [7:0] videosoc_csrbank12_tuning_word1_w;
wire videosoc_csrbank12_tuning_word0_re;
wire [7:0] videosoc_csrbank12_tuning_word0_r;
wire [7:0] videosoc_csrbank12_tuning_word0_w;
wire videosoc_csrbank12_sel;
reg comb_rhs_array_muxed0 = 1'd0;
reg [14:0] comb_rhs_array_muxed1 = 15'd0;
reg [2:0] comb_rhs_array_muxed2 = 3'd0;
reg comb_rhs_array_muxed3 = 1'd0;
reg comb_rhs_array_muxed4 = 1'd0;
reg comb_rhs_array_muxed5 = 1'd0;
reg comb_t_array_muxed0 = 1'd0;
reg comb_t_array_muxed1 = 1'd0;
reg comb_t_array_muxed2 = 1'd0;
reg comb_rhs_array_muxed6 = 1'd0;
reg [14:0] comb_rhs_array_muxed7 = 15'd0;
reg [2:0] comb_rhs_array_muxed8 = 3'd0;
reg comb_rhs_array_muxed9 = 1'd0;
reg comb_rhs_array_muxed10 = 1'd0;
reg comb_rhs_array_muxed11 = 1'd0;
reg comb_t_array_muxed3 = 1'd0;
reg comb_t_array_muxed4 = 1'd0;
reg comb_t_array_muxed5 = 1'd0;
reg [21:0] comb_rhs_array_muxed12 = 22'd0;
reg comb_rhs_array_muxed13 = 1'd0;
reg comb_rhs_array_muxed14 = 1'd0;
reg [21:0] comb_rhs_array_muxed15 = 22'd0;
reg comb_rhs_array_muxed16 = 1'd0;
reg comb_rhs_array_muxed17 = 1'd0;
reg [21:0] comb_rhs_array_muxed18 = 22'd0;
reg comb_rhs_array_muxed19 = 1'd0;
reg comb_rhs_array_muxed20 = 1'd0;
reg [21:0] comb_rhs_array_muxed21 = 22'd0;
reg comb_rhs_array_muxed22 = 1'd0;
reg comb_rhs_array_muxed23 = 1'd0;
reg [21:0] comb_rhs_array_muxed24 = 22'd0;
reg comb_rhs_array_muxed25 = 1'd0;
reg comb_rhs_array_muxed26 = 1'd0;
reg [21:0] comb_rhs_array_muxed27 = 22'd0;
reg comb_rhs_array_muxed28 = 1'd0;
reg comb_rhs_array_muxed29 = 1'd0;
reg [21:0] comb_rhs_array_muxed30 = 22'd0;
reg comb_rhs_array_muxed31 = 1'd0;
reg comb_rhs_array_muxed32 = 1'd0;
reg [21:0] comb_rhs_array_muxed33 = 22'd0;
reg comb_rhs_array_muxed34 = 1'd0;
reg comb_rhs_array_muxed35 = 1'd0;
reg [24:0] comb_rhs_array_muxed36 = 25'd0;
reg comb_rhs_array_muxed37 = 1'd0;
reg [29:0] comb_rhs_array_muxed38 = 30'd0;
reg [31:0] comb_rhs_array_muxed39 = 32'd0;
reg [3:0] comb_rhs_array_muxed40 = 4'd0;
reg comb_rhs_array_muxed41 = 1'd0;
reg comb_rhs_array_muxed42 = 1'd0;
reg comb_rhs_array_muxed43 = 1'd0;
reg [2:0] comb_rhs_array_muxed44 = 3'd0;
reg [1:0] comb_rhs_array_muxed45 = 2'd0;
reg [29:0] comb_rhs_array_muxed46 = 30'd0;
reg [31:0] comb_rhs_array_muxed47 = 32'd0;
reg [3:0] comb_rhs_array_muxed48 = 4'd0;
reg comb_rhs_array_muxed49 = 1'd0;
reg comb_rhs_array_muxed50 = 1'd0;
reg comb_rhs_array_muxed51 = 1'd0;
reg [2:0] comb_rhs_array_muxed52 = 3'd0;
reg [1:0] comb_rhs_array_muxed53 = 2'd0;
reg [9:0] sync_f_array_muxed0 = 10'd0;
reg [9:0] sync_f_array_muxed1 = 10'd0;
reg [9:0] sync_f_array_muxed2 = 10'd0;
reg [14:0] sync_rhs_array_muxed0 = 15'd0;
reg [2:0] sync_rhs_array_muxed1 = 3'd0;
reg sync_rhs_array_muxed2 = 1'd0;
reg sync_rhs_array_muxed3 = 1'd0;
reg sync_rhs_array_muxed4 = 1'd0;
reg sync_rhs_array_muxed5 = 1'd0;
reg sync_rhs_array_muxed6 = 1'd0;
reg [14:0] sync_rhs_array_muxed7 = 15'd0;
reg [2:0] sync_rhs_array_muxed8 = 3'd0;
reg sync_rhs_array_muxed9 = 1'd0;
reg sync_rhs_array_muxed10 = 1'd0;
reg sync_rhs_array_muxed11 = 1'd0;
reg sync_rhs_array_muxed12 = 1'd0;
reg sync_rhs_array_muxed13 = 1'd0;
reg [14:0] sync_rhs_array_muxed14 = 15'd0;
reg [2:0] sync_rhs_array_muxed15 = 3'd0;
reg sync_rhs_array_muxed16 = 1'd0;
reg sync_rhs_array_muxed17 = 1'd0;
reg sync_rhs_array_muxed18 = 1'd0;
reg sync_rhs_array_muxed19 = 1'd0;
reg sync_rhs_array_muxed20 = 1'd0;
reg [14:0] sync_rhs_array_muxed21 = 15'd0;
reg [2:0] sync_rhs_array_muxed22 = 3'd0;
reg sync_rhs_array_muxed23 = 1'd0;
reg sync_rhs_array_muxed24 = 1'd0;
reg sync_rhs_array_muxed25 = 1'd0;
reg sync_rhs_array_muxed26 = 1'd0;
reg sync_rhs_array_muxed27 = 1'd0;
(* ars_false_path = "true" *) wire xilinxasyncresetsynchronizerimpl0;
wire xilinxasyncresetsynchronizerimpl0_rst_meta;
(* ars_false_path = "true" *) wire xilinxasyncresetsynchronizerimpl1;
wire xilinxasyncresetsynchronizerimpl1_rst_meta;
(* ars_false_path = "true" *) wire xilinxasyncresetsynchronizerimpl2;
wire xilinxasyncresetsynchronizerimpl2_rst_meta;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl0_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl0_regs1 = 1'd0;
wire xilinxasyncresetsynchronizerimpl3_rst_meta;
wire xilinxasyncresetsynchronizerimpl4_rst_meta;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl1_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl1_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl2_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl2_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl3_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl3_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl4_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl4_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl5_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl5_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl6_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl6_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl7_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] xilinxmultiregimpl7_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl8_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl8_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl9_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl9_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl10_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl10_regs1 = 1'd0;
(* ars_false_path = "true" *) wire xilinxasyncresetsynchronizerimpl5;
wire xilinxasyncresetsynchronizerimpl5_rst_meta;
(* ars_false_path = "true" *) wire xilinxasyncresetsynchronizerimpl6;
wire xilinxasyncresetsynchronizerimpl6_rst_meta;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl11_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl11_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl12_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl12_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl13_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl13_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl14_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl14_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl15_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl15_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl16_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl16_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl17_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl17_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl18_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl18_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] xilinxmultiregimpl19_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] xilinxmultiregimpl19_regs1 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl20_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl20_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl21_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl21_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl22_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl22_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl23_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl23_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl24_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl24_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl25_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl25_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl26_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl26_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl27_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl27_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl28_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl28_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] xilinxmultiregimpl29_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] xilinxmultiregimpl29_regs1 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl30_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl30_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl31_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl31_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl32_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl32_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl33_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl33_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl34_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl34_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl35_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl35_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl36_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl36_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl37_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl37_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl38_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl38_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] xilinxmultiregimpl39_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] xilinxmultiregimpl39_regs1 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl40_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl40_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl41_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl41_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] xilinxmultiregimpl42_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] xilinxmultiregimpl42_regs1 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] xilinxmultiregimpl43_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] xilinxmultiregimpl43_regs1 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] xilinxmultiregimpl44_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] xilinxmultiregimpl44_regs1 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] xilinxmultiregimpl45_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] xilinxmultiregimpl45_regs1 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl46_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl46_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl47_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl47_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl48_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl48_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [5:0] xilinxmultiregimpl49_regs0 = 6'd0;
(* async_reg = "true", dont_touch = "true" *) reg [5:0] xilinxmultiregimpl49_regs1 = 6'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl50_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl50_regs1 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl51_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] xilinxmultiregimpl51_regs1 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] xilinxmultiregimpl52_regs0 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] xilinxmultiregimpl52_regs1 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] xilinxmultiregimpl53_regs0 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] xilinxmultiregimpl53_regs1 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl54_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl54_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl55_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] xilinxmultiregimpl55_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl56_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl56_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl57_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg xilinxmultiregimpl57_regs1 = 1'd0;

assign videosoc_sel = user_sw0;
assign hdmi_in0_freq_clk0 = hdmi_in0_pix_clk;
assign hdmi_in_txen = 1'd1;
always @(*) begin
	videosoc_videosoc_interrupt <= 32'd0;
	videosoc_videosoc_interrupt[1] <= videosoc_videosoc_irq;
	videosoc_videosoc_interrupt[2] <= videosoc_uart_irq;
	videosoc_videosoc_interrupt[3] <= ethmac_ev_irq;
	videosoc_videosoc_interrupt[4] <= dma_slot_array_irq;
end
assign videosoc_videosoc_ibus_adr = videosoc_videosoc_i_adr_o[31:2];
assign videosoc_videosoc_dbus_adr = videosoc_videosoc_d_adr_o[31:2];
assign videosoc_videosoc_rom_adr = videosoc_videosoc_rom_bus_adr[12:0];
assign videosoc_videosoc_rom_bus_dat_r = videosoc_videosoc_rom_dat_r;
always @(*) begin
	videosoc_videosoc_sram_we <= 4'd0;
	videosoc_videosoc_sram_we[0] <= (((videosoc_videosoc_sram_bus_cyc & videosoc_videosoc_sram_bus_stb) & videosoc_videosoc_sram_bus_we) & videosoc_videosoc_sram_bus_sel[0]);
	videosoc_videosoc_sram_we[1] <= (((videosoc_videosoc_sram_bus_cyc & videosoc_videosoc_sram_bus_stb) & videosoc_videosoc_sram_bus_we) & videosoc_videosoc_sram_bus_sel[1]);
	videosoc_videosoc_sram_we[2] <= (((videosoc_videosoc_sram_bus_cyc & videosoc_videosoc_sram_bus_stb) & videosoc_videosoc_sram_bus_we) & videosoc_videosoc_sram_bus_sel[2]);
	videosoc_videosoc_sram_we[3] <= (((videosoc_videosoc_sram_bus_cyc & videosoc_videosoc_sram_bus_stb) & videosoc_videosoc_sram_bus_we) & videosoc_videosoc_sram_bus_sel[3]);
end
assign videosoc_videosoc_sram_adr = videosoc_videosoc_sram_bus_adr[12:0];
assign videosoc_videosoc_sram_bus_dat_r = videosoc_videosoc_sram_dat_r;
assign videosoc_videosoc_sram_dat_w = videosoc_videosoc_sram_bus_dat_w;
assign videosoc_videosoc_zero_trigger = (videosoc_videosoc_value != 1'd0);
assign videosoc_videosoc_eventmanager_status_w = videosoc_videosoc_zero_status;
always @(*) begin
	videosoc_videosoc_zero_clear <= 1'd0;
	if ((videosoc_videosoc_eventmanager_pending_re & videosoc_videosoc_eventmanager_pending_r)) begin
		videosoc_videosoc_zero_clear <= 1'd1;
	end
end
assign videosoc_videosoc_eventmanager_pending_w = videosoc_videosoc_zero_pending;
assign videosoc_videosoc_irq = (videosoc_videosoc_eventmanager_pending_w & videosoc_videosoc_eventmanager_storage);
assign videosoc_videosoc_zero_status = videosoc_videosoc_zero_trigger;
assign videosoc_uart_tx_fifo_sink_valid = videosoc_uart_rxtx_re;
assign videosoc_uart_tx_fifo_sink_payload_data = videosoc_uart_rxtx_r;
assign videosoc_uart_txfull_status = (~videosoc_uart_tx_fifo_sink_ready);
assign videosoc_rs232phyinterface0_sink_valid = videosoc_uart_tx_fifo_source_valid;
assign videosoc_uart_tx_fifo_source_ready = videosoc_rs232phyinterface0_sink_ready;
assign videosoc_rs232phyinterface0_sink_first = videosoc_uart_tx_fifo_source_first;
assign videosoc_rs232phyinterface0_sink_last = videosoc_uart_tx_fifo_source_last;
assign videosoc_rs232phyinterface0_sink_payload_data = videosoc_uart_tx_fifo_source_payload_data;
assign videosoc_uart_tx_trigger = (~videosoc_uart_tx_fifo_sink_ready);
assign videosoc_uart_rx_fifo_sink_valid = videosoc_rs232phyinterface0_source_valid;
assign videosoc_rs232phyinterface0_source_ready = videosoc_uart_rx_fifo_sink_ready;
assign videosoc_uart_rx_fifo_sink_first = videosoc_rs232phyinterface0_source_first;
assign videosoc_uart_rx_fifo_sink_last = videosoc_rs232phyinterface0_source_last;
assign videosoc_uart_rx_fifo_sink_payload_data = videosoc_rs232phyinterface0_source_payload_data;
assign videosoc_uart_rxempty_status = (~videosoc_uart_rx_fifo_source_valid);
assign videosoc_uart_rxtx_w = videosoc_uart_rx_fifo_source_payload_data;
assign videosoc_uart_rx_fifo_source_ready = videosoc_uart_rx_clear;
assign videosoc_uart_rx_trigger = (~videosoc_uart_rx_fifo_source_valid);
always @(*) begin
	videosoc_uart_tx_clear <= 1'd0;
	if ((videosoc_uart_pending_re & videosoc_uart_pending_r[0])) begin
		videosoc_uart_tx_clear <= 1'd1;
	end
end
always @(*) begin
	videosoc_uart_status_w <= 2'd0;
	videosoc_uart_status_w[0] <= videosoc_uart_tx_status;
	videosoc_uart_status_w[1] <= videosoc_uart_rx_status;
end
always @(*) begin
	videosoc_uart_rx_clear <= 1'd0;
	if ((videosoc_uart_pending_re & videosoc_uart_pending_r[1])) begin
		videosoc_uart_rx_clear <= 1'd1;
	end
end
always @(*) begin
	videosoc_uart_pending_w <= 2'd0;
	videosoc_uart_pending_w[0] <= videosoc_uart_tx_pending;
	videosoc_uart_pending_w[1] <= videosoc_uart_rx_pending;
end
assign videosoc_uart_irq = ((videosoc_uart_pending_w[0] & videosoc_uart_storage[0]) | (videosoc_uart_pending_w[1] & videosoc_uart_storage[1]));
assign videosoc_uart_tx_status = videosoc_uart_tx_trigger;
assign videosoc_uart_rx_status = videosoc_uart_rx_trigger;
assign videosoc_uart_tx_fifo_syncfifo_din = {videosoc_uart_tx_fifo_fifo_in_last, videosoc_uart_tx_fifo_fifo_in_first, videosoc_uart_tx_fifo_fifo_in_payload_data};
assign {videosoc_uart_tx_fifo_fifo_out_last, videosoc_uart_tx_fifo_fifo_out_first, videosoc_uart_tx_fifo_fifo_out_payload_data} = videosoc_uart_tx_fifo_syncfifo_dout;
assign videosoc_uart_tx_fifo_sink_ready = videosoc_uart_tx_fifo_syncfifo_writable;
assign videosoc_uart_tx_fifo_syncfifo_we = videosoc_uart_tx_fifo_sink_valid;
assign videosoc_uart_tx_fifo_fifo_in_first = videosoc_uart_tx_fifo_sink_first;
assign videosoc_uart_tx_fifo_fifo_in_last = videosoc_uart_tx_fifo_sink_last;
assign videosoc_uart_tx_fifo_fifo_in_payload_data = videosoc_uart_tx_fifo_sink_payload_data;
assign videosoc_uart_tx_fifo_source_valid = videosoc_uart_tx_fifo_syncfifo_readable;
assign videosoc_uart_tx_fifo_source_first = videosoc_uart_tx_fifo_fifo_out_first;
assign videosoc_uart_tx_fifo_source_last = videosoc_uart_tx_fifo_fifo_out_last;
assign videosoc_uart_tx_fifo_source_payload_data = videosoc_uart_tx_fifo_fifo_out_payload_data;
assign videosoc_uart_tx_fifo_syncfifo_re = videosoc_uart_tx_fifo_source_ready;
always @(*) begin
	videosoc_uart_tx_fifo_wrport_adr <= 4'd0;
	if (videosoc_uart_tx_fifo_replace) begin
		videosoc_uart_tx_fifo_wrport_adr <= (videosoc_uart_tx_fifo_produce - 1'd1);
	end else begin
		videosoc_uart_tx_fifo_wrport_adr <= videosoc_uart_tx_fifo_produce;
	end
end
assign videosoc_uart_tx_fifo_wrport_dat_w = videosoc_uart_tx_fifo_syncfifo_din;
assign videosoc_uart_tx_fifo_wrport_we = (videosoc_uart_tx_fifo_syncfifo_we & (videosoc_uart_tx_fifo_syncfifo_writable | videosoc_uart_tx_fifo_replace));
assign videosoc_uart_tx_fifo_do_read = (videosoc_uart_tx_fifo_syncfifo_readable & videosoc_uart_tx_fifo_syncfifo_re);
assign videosoc_uart_tx_fifo_rdport_adr = videosoc_uart_tx_fifo_consume;
assign videosoc_uart_tx_fifo_syncfifo_dout = videosoc_uart_tx_fifo_rdport_dat_r;
assign videosoc_uart_tx_fifo_syncfifo_writable = (videosoc_uart_tx_fifo_level != 5'd16);
assign videosoc_uart_tx_fifo_syncfifo_readable = (videosoc_uart_tx_fifo_level != 1'd0);
assign videosoc_uart_rx_fifo_syncfifo_din = {videosoc_uart_rx_fifo_fifo_in_last, videosoc_uart_rx_fifo_fifo_in_first, videosoc_uart_rx_fifo_fifo_in_payload_data};
assign {videosoc_uart_rx_fifo_fifo_out_last, videosoc_uart_rx_fifo_fifo_out_first, videosoc_uart_rx_fifo_fifo_out_payload_data} = videosoc_uart_rx_fifo_syncfifo_dout;
assign videosoc_uart_rx_fifo_sink_ready = videosoc_uart_rx_fifo_syncfifo_writable;
assign videosoc_uart_rx_fifo_syncfifo_we = videosoc_uart_rx_fifo_sink_valid;
assign videosoc_uart_rx_fifo_fifo_in_first = videosoc_uart_rx_fifo_sink_first;
assign videosoc_uart_rx_fifo_fifo_in_last = videosoc_uart_rx_fifo_sink_last;
assign videosoc_uart_rx_fifo_fifo_in_payload_data = videosoc_uart_rx_fifo_sink_payload_data;
assign videosoc_uart_rx_fifo_source_valid = videosoc_uart_rx_fifo_syncfifo_readable;
assign videosoc_uart_rx_fifo_source_first = videosoc_uart_rx_fifo_fifo_out_first;
assign videosoc_uart_rx_fifo_source_last = videosoc_uart_rx_fifo_fifo_out_last;
assign videosoc_uart_rx_fifo_source_payload_data = videosoc_uart_rx_fifo_fifo_out_payload_data;
assign videosoc_uart_rx_fifo_syncfifo_re = videosoc_uart_rx_fifo_source_ready;
always @(*) begin
	videosoc_uart_rx_fifo_wrport_adr <= 4'd0;
	if (videosoc_uart_rx_fifo_replace) begin
		videosoc_uart_rx_fifo_wrport_adr <= (videosoc_uart_rx_fifo_produce - 1'd1);
	end else begin
		videosoc_uart_rx_fifo_wrport_adr <= videosoc_uart_rx_fifo_produce;
	end
end
assign videosoc_uart_rx_fifo_wrport_dat_w = videosoc_uart_rx_fifo_syncfifo_din;
assign videosoc_uart_rx_fifo_wrport_we = (videosoc_uart_rx_fifo_syncfifo_we & (videosoc_uart_rx_fifo_syncfifo_writable | videosoc_uart_rx_fifo_replace));
assign videosoc_uart_rx_fifo_do_read = (videosoc_uart_rx_fifo_syncfifo_readable & videosoc_uart_rx_fifo_syncfifo_re);
assign videosoc_uart_rx_fifo_rdport_adr = videosoc_uart_rx_fifo_consume;
assign videosoc_uart_rx_fifo_syncfifo_dout = videosoc_uart_rx_fifo_rdport_dat_r;
assign videosoc_uart_rx_fifo_syncfifo_writable = (videosoc_uart_rx_fifo_level != 5'd16);
assign videosoc_uart_rx_fifo_syncfifo_readable = (videosoc_uart_rx_fifo_level != 1'd0);
assign videosoc_bridge_reset = videosoc_bridge_done;
assign videosoc_rs232phyinterface1_source_ready = 1'd1;
assign videosoc_bridge_wishbone_adr = (videosoc_bridge_address + videosoc_bridge_word_counter);
assign videosoc_bridge_wishbone_dat_w = videosoc_bridge_data;
assign videosoc_bridge_wishbone_sel = 4'd15;
always @(*) begin
	videosoc_rs232phyinterface1_sink_payload_data <= 8'd0;
	case (videosoc_bridge_byte_counter)
		1'd0: begin
			videosoc_rs232phyinterface1_sink_payload_data <= videosoc_bridge_data[31:24];
		end
		1'd1: begin
			videosoc_rs232phyinterface1_sink_payload_data <= videosoc_bridge_data[23:16];
		end
		2'd2: begin
			videosoc_rs232phyinterface1_sink_payload_data <= videosoc_bridge_data[15:8];
		end
		default: begin
			videosoc_rs232phyinterface1_sink_payload_data <= videosoc_bridge_data[7:0];
		end
	endcase
end
assign videosoc_bridge_wait = (~videosoc_bridge_is_ongoing);
assign videosoc_rs232phyinterface1_sink_last = ((videosoc_bridge_byte_counter == 2'd3) & (videosoc_bridge_word_counter == (videosoc_bridge_length - 1'd1)));
always @(*) begin
	videosoc_bridge_wishbone_cyc <= 1'd0;
	videosoc_bridge_wishbone_stb <= 1'd0;
	videosoc_bridge_cmd_ce <= 1'd0;
	videosoc_bridge_is_ongoing <= 1'd0;
	videosoc_bridge_length_ce <= 1'd0;
	videosoc_bridge_wishbone_we <= 1'd0;
	videosoc_bridge_address_ce <= 1'd0;
	videosoc_bridge_word_counter_ce <= 1'd0;
	videosoc_rs232phyinterface1_sink_valid <= 1'd0;
	videosoc_bridge_rx_data_ce <= 1'd0;
	videosoc_bridge_byte_counter_reset <= 1'd0;
	videosoc_bridge_tx_data_ce <= 1'd0;
	videosoc_bridge_byte_counter_ce <= 1'd0;
	videosoc_bridge_word_counter_reset <= 1'd0;
	wishbonestreamingbridge_next_state <= 3'd0;
	wishbonestreamingbridge_next_state <= wishbonestreamingbridge_state;
	case (wishbonestreamingbridge_state)
		1'd1: begin
			if (videosoc_rs232phyinterface1_source_valid) begin
				videosoc_bridge_length_ce <= 1'd1;
				wishbonestreamingbridge_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (videosoc_rs232phyinterface1_source_valid) begin
				videosoc_bridge_address_ce <= 1'd1;
				videosoc_bridge_byte_counter_ce <= 1'd1;
				if ((videosoc_bridge_byte_counter == 2'd3)) begin
					if ((videosoc_bridge_cmd == 1'd1)) begin
						wishbonestreamingbridge_next_state <= 2'd3;
					end else begin
						if ((videosoc_bridge_cmd == 2'd2)) begin
							wishbonestreamingbridge_next_state <= 3'd5;
						end
					end
					videosoc_bridge_byte_counter_reset <= 1'd1;
				end
			end
		end
		2'd3: begin
			if (videosoc_rs232phyinterface1_source_valid) begin
				videosoc_bridge_rx_data_ce <= 1'd1;
				videosoc_bridge_byte_counter_ce <= 1'd1;
				if ((videosoc_bridge_byte_counter == 2'd3)) begin
					wishbonestreamingbridge_next_state <= 3'd4;
					videosoc_bridge_byte_counter_reset <= 1'd1;
				end
			end
		end
		3'd4: begin
			videosoc_bridge_wishbone_stb <= 1'd1;
			videosoc_bridge_wishbone_we <= 1'd1;
			videosoc_bridge_wishbone_cyc <= 1'd1;
			if (videosoc_bridge_wishbone_ack) begin
				videosoc_bridge_word_counter_ce <= 1'd1;
				if ((videosoc_bridge_word_counter == (videosoc_bridge_length - 1'd1))) begin
					wishbonestreamingbridge_next_state <= 1'd0;
				end else begin
					wishbonestreamingbridge_next_state <= 2'd3;
				end
			end
		end
		3'd5: begin
			videosoc_bridge_wishbone_stb <= 1'd1;
			videosoc_bridge_wishbone_we <= 1'd0;
			videosoc_bridge_wishbone_cyc <= 1'd1;
			if (videosoc_bridge_wishbone_ack) begin
				videosoc_bridge_tx_data_ce <= 1'd1;
				wishbonestreamingbridge_next_state <= 3'd6;
			end
		end
		3'd6: begin
			videosoc_rs232phyinterface1_sink_valid <= 1'd1;
			if (videosoc_rs232phyinterface1_sink_ready) begin
				videosoc_bridge_byte_counter_ce <= 1'd1;
				if ((videosoc_bridge_byte_counter == 2'd3)) begin
					videosoc_bridge_word_counter_ce <= 1'd1;
					if ((videosoc_bridge_word_counter == (videosoc_bridge_length - 1'd1))) begin
						wishbonestreamingbridge_next_state <= 1'd0;
					end else begin
						wishbonestreamingbridge_next_state <= 3'd5;
						videosoc_bridge_byte_counter_reset <= 1'd1;
					end
				end
			end
		end
		default: begin
			if (videosoc_rs232phyinterface1_source_valid) begin
				videosoc_bridge_cmd_ce <= 1'd1;
				if (((videosoc_rs232phyinterface1_source_payload_data == 1'd1) | (videosoc_rs232phyinterface1_source_payload_data == 2'd2))) begin
					wishbonestreamingbridge_next_state <= 1'd1;
				end
				videosoc_bridge_byte_counter_reset <= 1'd1;
				videosoc_bridge_word_counter_reset <= 1'd1;
			end
			videosoc_bridge_is_ongoing <= 1'd1;
		end
	endcase
end
assign videosoc_bridge_done = (videosoc_bridge_count == 1'd0);
always @(*) begin
	videosoc_rs232phyinterface0_source_valid <= 1'd0;
	videosoc_uart_phy_source_ready <= 1'd0;
	videosoc_rs232phyinterface0_source_first <= 1'd0;
	videosoc_rs232phyinterface0_source_last <= 1'd0;
	videosoc_rs232phyinterface0_source_payload_data <= 8'd0;
	videosoc_rs232phyinterface1_sink_ready <= 1'd0;
	videosoc_uart_phy_sink_valid <= 1'd0;
	videosoc_rs232phyinterface1_source_first <= 1'd0;
	videosoc_uart_phy_sink_first <= 1'd0;
	videosoc_rs232phyinterface1_source_valid <= 1'd0;
	videosoc_uart_phy_sink_last <= 1'd0;
	videosoc_uart_phy_sink_payload_data <= 8'd0;
	videosoc_rs232phyinterface0_sink_ready <= 1'd0;
	videosoc_rs232phyinterface1_source_last <= 1'd0;
	videosoc_rs232phyinterface1_source_payload_data <= 8'd0;
	videosoc_rs232phyinterface0_sink_ready <= 1'd1;
	videosoc_rs232phyinterface1_sink_ready <= 1'd1;
	case (videosoc_sel)
		1'd0: begin
			videosoc_rs232phyinterface0_source_valid <= videosoc_uart_phy_source_valid;
			videosoc_uart_phy_source_ready <= videosoc_rs232phyinterface0_source_ready;
			videosoc_rs232phyinterface0_source_first <= videosoc_uart_phy_source_first;
			videosoc_rs232phyinterface0_source_last <= videosoc_uart_phy_source_last;
			videosoc_rs232phyinterface0_source_payload_data <= videosoc_uart_phy_source_payload_data;
			videosoc_uart_phy_sink_valid <= videosoc_rs232phyinterface0_sink_valid;
			videosoc_rs232phyinterface0_sink_ready <= videosoc_uart_phy_sink_ready;
			videosoc_uart_phy_sink_first <= videosoc_rs232phyinterface0_sink_first;
			videosoc_uart_phy_sink_last <= videosoc_rs232phyinterface0_sink_last;
			videosoc_uart_phy_sink_payload_data <= videosoc_rs232phyinterface0_sink_payload_data;
		end
		1'd1: begin
			videosoc_rs232phyinterface1_source_valid <= videosoc_uart_phy_source_valid;
			videosoc_uart_phy_source_ready <= videosoc_rs232phyinterface1_source_ready;
			videosoc_rs232phyinterface1_source_first <= videosoc_uart_phy_source_first;
			videosoc_rs232phyinterface1_source_last <= videosoc_uart_phy_source_last;
			videosoc_rs232phyinterface1_source_payload_data <= videosoc_uart_phy_source_payload_data;
			videosoc_uart_phy_sink_valid <= videosoc_rs232phyinterface1_sink_valid;
			videosoc_rs232phyinterface1_sink_ready <= videosoc_uart_phy_sink_ready;
			videosoc_uart_phy_sink_first <= videosoc_rs232phyinterface1_sink_first;
			videosoc_uart_phy_sink_last <= videosoc_rs232phyinterface1_sink_last;
			videosoc_uart_phy_sink_payload_data <= videosoc_rs232phyinterface1_sink_payload_data;
		end
	endcase
end
assign videosoc_info_git_status = 160'd861173277431033699579123614235148681532316905970;
assign videosoc_info_platform_status = 63'd7954896779841861225;
assign videosoc_info_target_status = 63'd8532461355846860800;
assign oled_sclk = videosoc_oled_spi_pads_clk;
assign oled_sdin = videosoc_oled_spi_pads_mosi;
assign videosoc_oled_spimaster_start = (videosoc_oled_spimaster_ctrl_re & videosoc_oled_spimaster_ctrl_r);
assign videosoc_oled_spimaster_status = videosoc_oled_spimaster_done;
assign videosoc_oled_spimaster_set_clk = (videosoc_oled_spimaster_i == 3'd7);
assign videosoc_oled_spimaster_clr_clk = (videosoc_oled_spimaster_i == 4'd15);
assign videosoc_oled_spi_pads_cs_n = (~videosoc_oled_spimaster_enable_cs);
always @(*) begin
	videosoc_oled_spimaster_enable_shift <= 1'd0;
	oled_next_state <= 2'd0;
	videosoc_oled_spimaster_done <= 1'd0;
	videosoc_oled_spimaster_clr_cnt <= 1'd0;
	videosoc_oled_spimaster_inc_cnt <= 1'd0;
	videosoc_oled_spimaster_irq <= 1'd0;
	videosoc_oled_spimaster_enable_cs <= 1'd0;
	oled_next_state <= oled_state;
	case (oled_state)
		1'd1: begin
			if (videosoc_oled_spimaster_clr_clk) begin
				oled_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((videosoc_oled_spimaster_cnt == videosoc_oled_spimaster_length_storage)) begin
				oled_next_state <= 2'd3;
			end else begin
				videosoc_oled_spimaster_inc_cnt <= videosoc_oled_spimaster_clr_clk;
			end
			videosoc_oled_spimaster_enable_cs <= 1'd1;
			videosoc_oled_spimaster_enable_shift <= 1'd1;
		end
		2'd3: begin
			if (videosoc_oled_spimaster_set_clk) begin
				oled_next_state <= 1'd0;
			end
			videosoc_oled_spimaster_enable_shift <= 1'd1;
			videosoc_oled_spimaster_irq <= 1'd1;
		end
		default: begin
			if (videosoc_oled_spimaster_start) begin
				oled_next_state <= 1'd1;
			end
			videosoc_oled_spimaster_done <= 1'd1;
			videosoc_oled_spimaster_clr_cnt <= 1'd1;
		end
	endcase
end
assign {oled_vdd, oled_vbat, oled_dc, oled_res} = videosoc_oled_storage;
assign videosoc_ddrphy_oe = ((videosoc_ddrphy_last_wrdata_en[1] | videosoc_ddrphy_last_wrdata_en[2]) | videosoc_ddrphy_last_wrdata_en[3]);
assign videosoc_ddrphy_dfi_p0_address = videosoc_sdram_master_p0_address;
assign videosoc_ddrphy_dfi_p0_bank = videosoc_sdram_master_p0_bank;
assign videosoc_ddrphy_dfi_p0_cas_n = videosoc_sdram_master_p0_cas_n;
assign videosoc_ddrphy_dfi_p0_cs_n = videosoc_sdram_master_p0_cs_n;
assign videosoc_ddrphy_dfi_p0_ras_n = videosoc_sdram_master_p0_ras_n;
assign videosoc_ddrphy_dfi_p0_we_n = videosoc_sdram_master_p0_we_n;
assign videosoc_ddrphy_dfi_p0_cke = videosoc_sdram_master_p0_cke;
assign videosoc_ddrphy_dfi_p0_odt = videosoc_sdram_master_p0_odt;
assign videosoc_ddrphy_dfi_p0_reset_n = videosoc_sdram_master_p0_reset_n;
assign videosoc_ddrphy_dfi_p0_wrdata = videosoc_sdram_master_p0_wrdata;
assign videosoc_ddrphy_dfi_p0_wrdata_en = videosoc_sdram_master_p0_wrdata_en;
assign videosoc_ddrphy_dfi_p0_wrdata_mask = videosoc_sdram_master_p0_wrdata_mask;
assign videosoc_ddrphy_dfi_p0_rddata_en = videosoc_sdram_master_p0_rddata_en;
assign videosoc_sdram_master_p0_rddata = videosoc_ddrphy_dfi_p0_rddata;
assign videosoc_sdram_master_p0_rddata_valid = videosoc_ddrphy_dfi_p0_rddata_valid;
assign videosoc_ddrphy_dfi_p1_address = videosoc_sdram_master_p1_address;
assign videosoc_ddrphy_dfi_p1_bank = videosoc_sdram_master_p1_bank;
assign videosoc_ddrphy_dfi_p1_cas_n = videosoc_sdram_master_p1_cas_n;
assign videosoc_ddrphy_dfi_p1_cs_n = videosoc_sdram_master_p1_cs_n;
assign videosoc_ddrphy_dfi_p1_ras_n = videosoc_sdram_master_p1_ras_n;
assign videosoc_ddrphy_dfi_p1_we_n = videosoc_sdram_master_p1_we_n;
assign videosoc_ddrphy_dfi_p1_cke = videosoc_sdram_master_p1_cke;
assign videosoc_ddrphy_dfi_p1_odt = videosoc_sdram_master_p1_odt;
assign videosoc_ddrphy_dfi_p1_reset_n = videosoc_sdram_master_p1_reset_n;
assign videosoc_ddrphy_dfi_p1_wrdata = videosoc_sdram_master_p1_wrdata;
assign videosoc_ddrphy_dfi_p1_wrdata_en = videosoc_sdram_master_p1_wrdata_en;
assign videosoc_ddrphy_dfi_p1_wrdata_mask = videosoc_sdram_master_p1_wrdata_mask;
assign videosoc_ddrphy_dfi_p1_rddata_en = videosoc_sdram_master_p1_rddata_en;
assign videosoc_sdram_master_p1_rddata = videosoc_ddrphy_dfi_p1_rddata;
assign videosoc_sdram_master_p1_rddata_valid = videosoc_ddrphy_dfi_p1_rddata_valid;
assign videosoc_ddrphy_dfi_p2_address = videosoc_sdram_master_p2_address;
assign videosoc_ddrphy_dfi_p2_bank = videosoc_sdram_master_p2_bank;
assign videosoc_ddrphy_dfi_p2_cas_n = videosoc_sdram_master_p2_cas_n;
assign videosoc_ddrphy_dfi_p2_cs_n = videosoc_sdram_master_p2_cs_n;
assign videosoc_ddrphy_dfi_p2_ras_n = videosoc_sdram_master_p2_ras_n;
assign videosoc_ddrphy_dfi_p2_we_n = videosoc_sdram_master_p2_we_n;
assign videosoc_ddrphy_dfi_p2_cke = videosoc_sdram_master_p2_cke;
assign videosoc_ddrphy_dfi_p2_odt = videosoc_sdram_master_p2_odt;
assign videosoc_ddrphy_dfi_p2_reset_n = videosoc_sdram_master_p2_reset_n;
assign videosoc_ddrphy_dfi_p2_wrdata = videosoc_sdram_master_p2_wrdata;
assign videosoc_ddrphy_dfi_p2_wrdata_en = videosoc_sdram_master_p2_wrdata_en;
assign videosoc_ddrphy_dfi_p2_wrdata_mask = videosoc_sdram_master_p2_wrdata_mask;
assign videosoc_ddrphy_dfi_p2_rddata_en = videosoc_sdram_master_p2_rddata_en;
assign videosoc_sdram_master_p2_rddata = videosoc_ddrphy_dfi_p2_rddata;
assign videosoc_sdram_master_p2_rddata_valid = videosoc_ddrphy_dfi_p2_rddata_valid;
assign videosoc_ddrphy_dfi_p3_address = videosoc_sdram_master_p3_address;
assign videosoc_ddrphy_dfi_p3_bank = videosoc_sdram_master_p3_bank;
assign videosoc_ddrphy_dfi_p3_cas_n = videosoc_sdram_master_p3_cas_n;
assign videosoc_ddrphy_dfi_p3_cs_n = videosoc_sdram_master_p3_cs_n;
assign videosoc_ddrphy_dfi_p3_ras_n = videosoc_sdram_master_p3_ras_n;
assign videosoc_ddrphy_dfi_p3_we_n = videosoc_sdram_master_p3_we_n;
assign videosoc_ddrphy_dfi_p3_cke = videosoc_sdram_master_p3_cke;
assign videosoc_ddrphy_dfi_p3_odt = videosoc_sdram_master_p3_odt;
assign videosoc_ddrphy_dfi_p3_reset_n = videosoc_sdram_master_p3_reset_n;
assign videosoc_ddrphy_dfi_p3_wrdata = videosoc_sdram_master_p3_wrdata;
assign videosoc_ddrphy_dfi_p3_wrdata_en = videosoc_sdram_master_p3_wrdata_en;
assign videosoc_ddrphy_dfi_p3_wrdata_mask = videosoc_sdram_master_p3_wrdata_mask;
assign videosoc_ddrphy_dfi_p3_rddata_en = videosoc_sdram_master_p3_rddata_en;
assign videosoc_sdram_master_p3_rddata = videosoc_ddrphy_dfi_p3_rddata;
assign videosoc_sdram_master_p3_rddata_valid = videosoc_ddrphy_dfi_p3_rddata_valid;
assign videosoc_sdram_slave_p0_address = videosoc_sdram_dfi_p0_address;
assign videosoc_sdram_slave_p0_bank = videosoc_sdram_dfi_p0_bank;
assign videosoc_sdram_slave_p0_cas_n = videosoc_sdram_dfi_p0_cas_n;
assign videosoc_sdram_slave_p0_cs_n = videosoc_sdram_dfi_p0_cs_n;
assign videosoc_sdram_slave_p0_ras_n = videosoc_sdram_dfi_p0_ras_n;
assign videosoc_sdram_slave_p0_we_n = videosoc_sdram_dfi_p0_we_n;
assign videosoc_sdram_slave_p0_cke = videosoc_sdram_dfi_p0_cke;
assign videosoc_sdram_slave_p0_odt = videosoc_sdram_dfi_p0_odt;
assign videosoc_sdram_slave_p0_reset_n = videosoc_sdram_dfi_p0_reset_n;
assign videosoc_sdram_slave_p0_wrdata = videosoc_sdram_dfi_p0_wrdata;
assign videosoc_sdram_slave_p0_wrdata_en = videosoc_sdram_dfi_p0_wrdata_en;
assign videosoc_sdram_slave_p0_wrdata_mask = videosoc_sdram_dfi_p0_wrdata_mask;
assign videosoc_sdram_slave_p0_rddata_en = videosoc_sdram_dfi_p0_rddata_en;
assign videosoc_sdram_dfi_p0_rddata = videosoc_sdram_slave_p0_rddata;
assign videosoc_sdram_dfi_p0_rddata_valid = videosoc_sdram_slave_p0_rddata_valid;
assign videosoc_sdram_slave_p1_address = videosoc_sdram_dfi_p1_address;
assign videosoc_sdram_slave_p1_bank = videosoc_sdram_dfi_p1_bank;
assign videosoc_sdram_slave_p1_cas_n = videosoc_sdram_dfi_p1_cas_n;
assign videosoc_sdram_slave_p1_cs_n = videosoc_sdram_dfi_p1_cs_n;
assign videosoc_sdram_slave_p1_ras_n = videosoc_sdram_dfi_p1_ras_n;
assign videosoc_sdram_slave_p1_we_n = videosoc_sdram_dfi_p1_we_n;
assign videosoc_sdram_slave_p1_cke = videosoc_sdram_dfi_p1_cke;
assign videosoc_sdram_slave_p1_odt = videosoc_sdram_dfi_p1_odt;
assign videosoc_sdram_slave_p1_reset_n = videosoc_sdram_dfi_p1_reset_n;
assign videosoc_sdram_slave_p1_wrdata = videosoc_sdram_dfi_p1_wrdata;
assign videosoc_sdram_slave_p1_wrdata_en = videosoc_sdram_dfi_p1_wrdata_en;
assign videosoc_sdram_slave_p1_wrdata_mask = videosoc_sdram_dfi_p1_wrdata_mask;
assign videosoc_sdram_slave_p1_rddata_en = videosoc_sdram_dfi_p1_rddata_en;
assign videosoc_sdram_dfi_p1_rddata = videosoc_sdram_slave_p1_rddata;
assign videosoc_sdram_dfi_p1_rddata_valid = videosoc_sdram_slave_p1_rddata_valid;
assign videosoc_sdram_slave_p2_address = videosoc_sdram_dfi_p2_address;
assign videosoc_sdram_slave_p2_bank = videosoc_sdram_dfi_p2_bank;
assign videosoc_sdram_slave_p2_cas_n = videosoc_sdram_dfi_p2_cas_n;
assign videosoc_sdram_slave_p2_cs_n = videosoc_sdram_dfi_p2_cs_n;
assign videosoc_sdram_slave_p2_ras_n = videosoc_sdram_dfi_p2_ras_n;
assign videosoc_sdram_slave_p2_we_n = videosoc_sdram_dfi_p2_we_n;
assign videosoc_sdram_slave_p2_cke = videosoc_sdram_dfi_p2_cke;
assign videosoc_sdram_slave_p2_odt = videosoc_sdram_dfi_p2_odt;
assign videosoc_sdram_slave_p2_reset_n = videosoc_sdram_dfi_p2_reset_n;
assign videosoc_sdram_slave_p2_wrdata = videosoc_sdram_dfi_p2_wrdata;
assign videosoc_sdram_slave_p2_wrdata_en = videosoc_sdram_dfi_p2_wrdata_en;
assign videosoc_sdram_slave_p2_wrdata_mask = videosoc_sdram_dfi_p2_wrdata_mask;
assign videosoc_sdram_slave_p2_rddata_en = videosoc_sdram_dfi_p2_rddata_en;
assign videosoc_sdram_dfi_p2_rddata = videosoc_sdram_slave_p2_rddata;
assign videosoc_sdram_dfi_p2_rddata_valid = videosoc_sdram_slave_p2_rddata_valid;
assign videosoc_sdram_slave_p3_address = videosoc_sdram_dfi_p3_address;
assign videosoc_sdram_slave_p3_bank = videosoc_sdram_dfi_p3_bank;
assign videosoc_sdram_slave_p3_cas_n = videosoc_sdram_dfi_p3_cas_n;
assign videosoc_sdram_slave_p3_cs_n = videosoc_sdram_dfi_p3_cs_n;
assign videosoc_sdram_slave_p3_ras_n = videosoc_sdram_dfi_p3_ras_n;
assign videosoc_sdram_slave_p3_we_n = videosoc_sdram_dfi_p3_we_n;
assign videosoc_sdram_slave_p3_cke = videosoc_sdram_dfi_p3_cke;
assign videosoc_sdram_slave_p3_odt = videosoc_sdram_dfi_p3_odt;
assign videosoc_sdram_slave_p3_reset_n = videosoc_sdram_dfi_p3_reset_n;
assign videosoc_sdram_slave_p3_wrdata = videosoc_sdram_dfi_p3_wrdata;
assign videosoc_sdram_slave_p3_wrdata_en = videosoc_sdram_dfi_p3_wrdata_en;
assign videosoc_sdram_slave_p3_wrdata_mask = videosoc_sdram_dfi_p3_wrdata_mask;
assign videosoc_sdram_slave_p3_rddata_en = videosoc_sdram_dfi_p3_rddata_en;
assign videosoc_sdram_dfi_p3_rddata = videosoc_sdram_slave_p3_rddata;
assign videosoc_sdram_dfi_p3_rddata_valid = videosoc_sdram_slave_p3_rddata_valid;
always @(*) begin
	videosoc_sdram_master_p2_cs_n <= 1'd1;
	videosoc_sdram_master_p2_ras_n <= 1'd1;
	videosoc_sdram_master_p2_we_n <= 1'd1;
	videosoc_sdram_inti_p2_rddata <= 32'd0;
	videosoc_sdram_master_p2_cke <= 1'd0;
	videosoc_sdram_inti_p2_rddata_valid <= 1'd0;
	videosoc_sdram_master_p2_odt <= 1'd0;
	videosoc_sdram_master_p2_reset_n <= 1'd0;
	videosoc_sdram_master_p2_wrdata <= 32'd0;
	videosoc_sdram_master_p2_wrdata_en <= 1'd0;
	videosoc_sdram_master_p2_wrdata_mask <= 4'd0;
	videosoc_sdram_master_p2_rddata_en <= 1'd0;
	videosoc_sdram_master_p3_address <= 15'd0;
	videosoc_sdram_master_p3_bank <= 3'd0;
	videosoc_sdram_master_p3_cas_n <= 1'd1;
	videosoc_sdram_master_p3_cs_n <= 1'd1;
	videosoc_sdram_master_p3_ras_n <= 1'd1;
	videosoc_sdram_master_p3_we_n <= 1'd1;
	videosoc_sdram_inti_p3_rddata <= 32'd0;
	videosoc_sdram_master_p3_cke <= 1'd0;
	videosoc_sdram_inti_p3_rddata_valid <= 1'd0;
	videosoc_sdram_master_p3_odt <= 1'd0;
	videosoc_sdram_master_p3_reset_n <= 1'd0;
	videosoc_sdram_master_p3_wrdata <= 32'd0;
	videosoc_sdram_master_p3_wrdata_en <= 1'd0;
	videosoc_sdram_master_p3_wrdata_mask <= 4'd0;
	videosoc_sdram_master_p3_rddata_en <= 1'd0;
	videosoc_sdram_slave_p0_rddata <= 32'd0;
	videosoc_sdram_slave_p0_rddata_valid <= 1'd0;
	videosoc_sdram_slave_p1_rddata <= 32'd0;
	videosoc_sdram_slave_p1_rddata_valid <= 1'd0;
	videosoc_sdram_slave_p2_rddata <= 32'd0;
	videosoc_sdram_slave_p2_rddata_valid <= 1'd0;
	videosoc_sdram_slave_p3_rddata <= 32'd0;
	videosoc_sdram_slave_p3_rddata_valid <= 1'd0;
	videosoc_sdram_master_p0_address <= 15'd0;
	videosoc_sdram_master_p0_bank <= 3'd0;
	videosoc_sdram_master_p0_cas_n <= 1'd1;
	videosoc_sdram_master_p0_cs_n <= 1'd1;
	videosoc_sdram_master_p0_ras_n <= 1'd1;
	videosoc_sdram_master_p0_we_n <= 1'd1;
	videosoc_sdram_inti_p0_rddata <= 32'd0;
	videosoc_sdram_master_p0_cke <= 1'd0;
	videosoc_sdram_inti_p0_rddata_valid <= 1'd0;
	videosoc_sdram_master_p0_odt <= 1'd0;
	videosoc_sdram_master_p0_reset_n <= 1'd0;
	videosoc_sdram_master_p0_wrdata <= 32'd0;
	videosoc_sdram_master_p0_wrdata_en <= 1'd0;
	videosoc_sdram_master_p0_wrdata_mask <= 4'd0;
	videosoc_sdram_master_p0_rddata_en <= 1'd0;
	videosoc_sdram_master_p1_address <= 15'd0;
	videosoc_sdram_master_p1_bank <= 3'd0;
	videosoc_sdram_master_p1_cas_n <= 1'd1;
	videosoc_sdram_master_p1_cs_n <= 1'd1;
	videosoc_sdram_master_p1_ras_n <= 1'd1;
	videosoc_sdram_master_p1_we_n <= 1'd1;
	videosoc_sdram_inti_p1_rddata <= 32'd0;
	videosoc_sdram_master_p1_cke <= 1'd0;
	videosoc_sdram_inti_p1_rddata_valid <= 1'd0;
	videosoc_sdram_master_p1_odt <= 1'd0;
	videosoc_sdram_master_p1_reset_n <= 1'd0;
	videosoc_sdram_master_p1_wrdata <= 32'd0;
	videosoc_sdram_master_p1_wrdata_en <= 1'd0;
	videosoc_sdram_master_p1_wrdata_mask <= 4'd0;
	videosoc_sdram_master_p1_rddata_en <= 1'd0;
	videosoc_sdram_master_p2_address <= 15'd0;
	videosoc_sdram_master_p2_bank <= 3'd0;
	videosoc_sdram_master_p2_cas_n <= 1'd1;
	if (videosoc_sdram_storage[0]) begin
		videosoc_sdram_master_p0_address <= videosoc_sdram_slave_p0_address;
		videosoc_sdram_master_p0_bank <= videosoc_sdram_slave_p0_bank;
		videosoc_sdram_master_p0_cas_n <= videosoc_sdram_slave_p0_cas_n;
		videosoc_sdram_master_p0_cs_n <= videosoc_sdram_slave_p0_cs_n;
		videosoc_sdram_master_p0_ras_n <= videosoc_sdram_slave_p0_ras_n;
		videosoc_sdram_master_p0_we_n <= videosoc_sdram_slave_p0_we_n;
		videosoc_sdram_master_p0_cke <= videosoc_sdram_slave_p0_cke;
		videosoc_sdram_master_p0_odt <= videosoc_sdram_slave_p0_odt;
		videosoc_sdram_master_p0_reset_n <= videosoc_sdram_slave_p0_reset_n;
		videosoc_sdram_master_p0_wrdata <= videosoc_sdram_slave_p0_wrdata;
		videosoc_sdram_master_p0_wrdata_en <= videosoc_sdram_slave_p0_wrdata_en;
		videosoc_sdram_master_p0_wrdata_mask <= videosoc_sdram_slave_p0_wrdata_mask;
		videosoc_sdram_master_p0_rddata_en <= videosoc_sdram_slave_p0_rddata_en;
		videosoc_sdram_slave_p0_rddata <= videosoc_sdram_master_p0_rddata;
		videosoc_sdram_slave_p0_rddata_valid <= videosoc_sdram_master_p0_rddata_valid;
		videosoc_sdram_master_p1_address <= videosoc_sdram_slave_p1_address;
		videosoc_sdram_master_p1_bank <= videosoc_sdram_slave_p1_bank;
		videosoc_sdram_master_p1_cas_n <= videosoc_sdram_slave_p1_cas_n;
		videosoc_sdram_master_p1_cs_n <= videosoc_sdram_slave_p1_cs_n;
		videosoc_sdram_master_p1_ras_n <= videosoc_sdram_slave_p1_ras_n;
		videosoc_sdram_master_p1_we_n <= videosoc_sdram_slave_p1_we_n;
		videosoc_sdram_master_p1_cke <= videosoc_sdram_slave_p1_cke;
		videosoc_sdram_master_p1_odt <= videosoc_sdram_slave_p1_odt;
		videosoc_sdram_master_p1_reset_n <= videosoc_sdram_slave_p1_reset_n;
		videosoc_sdram_master_p1_wrdata <= videosoc_sdram_slave_p1_wrdata;
		videosoc_sdram_master_p1_wrdata_en <= videosoc_sdram_slave_p1_wrdata_en;
		videosoc_sdram_master_p1_wrdata_mask <= videosoc_sdram_slave_p1_wrdata_mask;
		videosoc_sdram_master_p1_rddata_en <= videosoc_sdram_slave_p1_rddata_en;
		videosoc_sdram_slave_p1_rddata <= videosoc_sdram_master_p1_rddata;
		videosoc_sdram_slave_p1_rddata_valid <= videosoc_sdram_master_p1_rddata_valid;
		videosoc_sdram_master_p2_address <= videosoc_sdram_slave_p2_address;
		videosoc_sdram_master_p2_bank <= videosoc_sdram_slave_p2_bank;
		videosoc_sdram_master_p2_cas_n <= videosoc_sdram_slave_p2_cas_n;
		videosoc_sdram_master_p2_cs_n <= videosoc_sdram_slave_p2_cs_n;
		videosoc_sdram_master_p2_ras_n <= videosoc_sdram_slave_p2_ras_n;
		videosoc_sdram_master_p2_we_n <= videosoc_sdram_slave_p2_we_n;
		videosoc_sdram_master_p2_cke <= videosoc_sdram_slave_p2_cke;
		videosoc_sdram_master_p2_odt <= videosoc_sdram_slave_p2_odt;
		videosoc_sdram_master_p2_reset_n <= videosoc_sdram_slave_p2_reset_n;
		videosoc_sdram_master_p2_wrdata <= videosoc_sdram_slave_p2_wrdata;
		videosoc_sdram_master_p2_wrdata_en <= videosoc_sdram_slave_p2_wrdata_en;
		videosoc_sdram_master_p2_wrdata_mask <= videosoc_sdram_slave_p2_wrdata_mask;
		videosoc_sdram_master_p2_rddata_en <= videosoc_sdram_slave_p2_rddata_en;
		videosoc_sdram_slave_p2_rddata <= videosoc_sdram_master_p2_rddata;
		videosoc_sdram_slave_p2_rddata_valid <= videosoc_sdram_master_p2_rddata_valid;
		videosoc_sdram_master_p3_address <= videosoc_sdram_slave_p3_address;
		videosoc_sdram_master_p3_bank <= videosoc_sdram_slave_p3_bank;
		videosoc_sdram_master_p3_cas_n <= videosoc_sdram_slave_p3_cas_n;
		videosoc_sdram_master_p3_cs_n <= videosoc_sdram_slave_p3_cs_n;
		videosoc_sdram_master_p3_ras_n <= videosoc_sdram_slave_p3_ras_n;
		videosoc_sdram_master_p3_we_n <= videosoc_sdram_slave_p3_we_n;
		videosoc_sdram_master_p3_cke <= videosoc_sdram_slave_p3_cke;
		videosoc_sdram_master_p3_odt <= videosoc_sdram_slave_p3_odt;
		videosoc_sdram_master_p3_reset_n <= videosoc_sdram_slave_p3_reset_n;
		videosoc_sdram_master_p3_wrdata <= videosoc_sdram_slave_p3_wrdata;
		videosoc_sdram_master_p3_wrdata_en <= videosoc_sdram_slave_p3_wrdata_en;
		videosoc_sdram_master_p3_wrdata_mask <= videosoc_sdram_slave_p3_wrdata_mask;
		videosoc_sdram_master_p3_rddata_en <= videosoc_sdram_slave_p3_rddata_en;
		videosoc_sdram_slave_p3_rddata <= videosoc_sdram_master_p3_rddata;
		videosoc_sdram_slave_p3_rddata_valid <= videosoc_sdram_master_p3_rddata_valid;
	end else begin
		videosoc_sdram_master_p0_address <= videosoc_sdram_inti_p0_address;
		videosoc_sdram_master_p0_bank <= videosoc_sdram_inti_p0_bank;
		videosoc_sdram_master_p0_cas_n <= videosoc_sdram_inti_p0_cas_n;
		videosoc_sdram_master_p0_cs_n <= videosoc_sdram_inti_p0_cs_n;
		videosoc_sdram_master_p0_ras_n <= videosoc_sdram_inti_p0_ras_n;
		videosoc_sdram_master_p0_we_n <= videosoc_sdram_inti_p0_we_n;
		videosoc_sdram_master_p0_cke <= videosoc_sdram_inti_p0_cke;
		videosoc_sdram_master_p0_odt <= videosoc_sdram_inti_p0_odt;
		videosoc_sdram_master_p0_reset_n <= videosoc_sdram_inti_p0_reset_n;
		videosoc_sdram_master_p0_wrdata <= videosoc_sdram_inti_p0_wrdata;
		videosoc_sdram_master_p0_wrdata_en <= videosoc_sdram_inti_p0_wrdata_en;
		videosoc_sdram_master_p0_wrdata_mask <= videosoc_sdram_inti_p0_wrdata_mask;
		videosoc_sdram_master_p0_rddata_en <= videosoc_sdram_inti_p0_rddata_en;
		videosoc_sdram_inti_p0_rddata <= videosoc_sdram_master_p0_rddata;
		videosoc_sdram_inti_p0_rddata_valid <= videosoc_sdram_master_p0_rddata_valid;
		videosoc_sdram_master_p1_address <= videosoc_sdram_inti_p1_address;
		videosoc_sdram_master_p1_bank <= videosoc_sdram_inti_p1_bank;
		videosoc_sdram_master_p1_cas_n <= videosoc_sdram_inti_p1_cas_n;
		videosoc_sdram_master_p1_cs_n <= videosoc_sdram_inti_p1_cs_n;
		videosoc_sdram_master_p1_ras_n <= videosoc_sdram_inti_p1_ras_n;
		videosoc_sdram_master_p1_we_n <= videosoc_sdram_inti_p1_we_n;
		videosoc_sdram_master_p1_cke <= videosoc_sdram_inti_p1_cke;
		videosoc_sdram_master_p1_odt <= videosoc_sdram_inti_p1_odt;
		videosoc_sdram_master_p1_reset_n <= videosoc_sdram_inti_p1_reset_n;
		videosoc_sdram_master_p1_wrdata <= videosoc_sdram_inti_p1_wrdata;
		videosoc_sdram_master_p1_wrdata_en <= videosoc_sdram_inti_p1_wrdata_en;
		videosoc_sdram_master_p1_wrdata_mask <= videosoc_sdram_inti_p1_wrdata_mask;
		videosoc_sdram_master_p1_rddata_en <= videosoc_sdram_inti_p1_rddata_en;
		videosoc_sdram_inti_p1_rddata <= videosoc_sdram_master_p1_rddata;
		videosoc_sdram_inti_p1_rddata_valid <= videosoc_sdram_master_p1_rddata_valid;
		videosoc_sdram_master_p2_address <= videosoc_sdram_inti_p2_address;
		videosoc_sdram_master_p2_bank <= videosoc_sdram_inti_p2_bank;
		videosoc_sdram_master_p2_cas_n <= videosoc_sdram_inti_p2_cas_n;
		videosoc_sdram_master_p2_cs_n <= videosoc_sdram_inti_p2_cs_n;
		videosoc_sdram_master_p2_ras_n <= videosoc_sdram_inti_p2_ras_n;
		videosoc_sdram_master_p2_we_n <= videosoc_sdram_inti_p2_we_n;
		videosoc_sdram_master_p2_cke <= videosoc_sdram_inti_p2_cke;
		videosoc_sdram_master_p2_odt <= videosoc_sdram_inti_p2_odt;
		videosoc_sdram_master_p2_reset_n <= videosoc_sdram_inti_p2_reset_n;
		videosoc_sdram_master_p2_wrdata <= videosoc_sdram_inti_p2_wrdata;
		videosoc_sdram_master_p2_wrdata_en <= videosoc_sdram_inti_p2_wrdata_en;
		videosoc_sdram_master_p2_wrdata_mask <= videosoc_sdram_inti_p2_wrdata_mask;
		videosoc_sdram_master_p2_rddata_en <= videosoc_sdram_inti_p2_rddata_en;
		videosoc_sdram_inti_p2_rddata <= videosoc_sdram_master_p2_rddata;
		videosoc_sdram_inti_p2_rddata_valid <= videosoc_sdram_master_p2_rddata_valid;
		videosoc_sdram_master_p3_address <= videosoc_sdram_inti_p3_address;
		videosoc_sdram_master_p3_bank <= videosoc_sdram_inti_p3_bank;
		videosoc_sdram_master_p3_cas_n <= videosoc_sdram_inti_p3_cas_n;
		videosoc_sdram_master_p3_cs_n <= videosoc_sdram_inti_p3_cs_n;
		videosoc_sdram_master_p3_ras_n <= videosoc_sdram_inti_p3_ras_n;
		videosoc_sdram_master_p3_we_n <= videosoc_sdram_inti_p3_we_n;
		videosoc_sdram_master_p3_cke <= videosoc_sdram_inti_p3_cke;
		videosoc_sdram_master_p3_odt <= videosoc_sdram_inti_p3_odt;
		videosoc_sdram_master_p3_reset_n <= videosoc_sdram_inti_p3_reset_n;
		videosoc_sdram_master_p3_wrdata <= videosoc_sdram_inti_p3_wrdata;
		videosoc_sdram_master_p3_wrdata_en <= videosoc_sdram_inti_p3_wrdata_en;
		videosoc_sdram_master_p3_wrdata_mask <= videosoc_sdram_inti_p3_wrdata_mask;
		videosoc_sdram_master_p3_rddata_en <= videosoc_sdram_inti_p3_rddata_en;
		videosoc_sdram_inti_p3_rddata <= videosoc_sdram_master_p3_rddata;
		videosoc_sdram_inti_p3_rddata_valid <= videosoc_sdram_master_p3_rddata_valid;
	end
end
assign videosoc_sdram_inti_p0_cke = videosoc_sdram_storage[1];
assign videosoc_sdram_inti_p1_cke = videosoc_sdram_storage[1];
assign videosoc_sdram_inti_p2_cke = videosoc_sdram_storage[1];
assign videosoc_sdram_inti_p3_cke = videosoc_sdram_storage[1];
assign videosoc_sdram_inti_p0_odt = videosoc_sdram_storage[2];
assign videosoc_sdram_inti_p1_odt = videosoc_sdram_storage[2];
assign videosoc_sdram_inti_p2_odt = videosoc_sdram_storage[2];
assign videosoc_sdram_inti_p3_odt = videosoc_sdram_storage[2];
assign videosoc_sdram_inti_p0_reset_n = videosoc_sdram_storage[3];
assign videosoc_sdram_inti_p1_reset_n = videosoc_sdram_storage[3];
assign videosoc_sdram_inti_p2_reset_n = videosoc_sdram_storage[3];
assign videosoc_sdram_inti_p3_reset_n = videosoc_sdram_storage[3];
always @(*) begin
	videosoc_sdram_inti_p0_we_n <= 1'd1;
	videosoc_sdram_inti_p0_cas_n <= 1'd1;
	videosoc_sdram_inti_p0_cs_n <= 1'd1;
	videosoc_sdram_inti_p0_ras_n <= 1'd1;
	if (videosoc_sdram_phaseinjector0_command_issue_re) begin
		videosoc_sdram_inti_p0_cs_n <= (~videosoc_sdram_phaseinjector0_command_storage[0]);
		videosoc_sdram_inti_p0_we_n <= (~videosoc_sdram_phaseinjector0_command_storage[1]);
		videosoc_sdram_inti_p0_cas_n <= (~videosoc_sdram_phaseinjector0_command_storage[2]);
		videosoc_sdram_inti_p0_ras_n <= (~videosoc_sdram_phaseinjector0_command_storage[3]);
	end else begin
		videosoc_sdram_inti_p0_cs_n <= 1'd1;
		videosoc_sdram_inti_p0_we_n <= 1'd1;
		videosoc_sdram_inti_p0_cas_n <= 1'd1;
		videosoc_sdram_inti_p0_ras_n <= 1'd1;
	end
end
assign videosoc_sdram_inti_p0_address = videosoc_sdram_phaseinjector0_address_storage;
assign videosoc_sdram_inti_p0_bank = videosoc_sdram_phaseinjector0_baddress_storage;
assign videosoc_sdram_inti_p0_wrdata_en = (videosoc_sdram_phaseinjector0_command_issue_re & videosoc_sdram_phaseinjector0_command_storage[4]);
assign videosoc_sdram_inti_p0_rddata_en = (videosoc_sdram_phaseinjector0_command_issue_re & videosoc_sdram_phaseinjector0_command_storage[5]);
assign videosoc_sdram_inti_p0_wrdata = videosoc_sdram_phaseinjector0_wrdata_storage;
assign videosoc_sdram_inti_p0_wrdata_mask = 1'd0;
always @(*) begin
	videosoc_sdram_inti_p1_cas_n <= 1'd1;
	videosoc_sdram_inti_p1_cs_n <= 1'd1;
	videosoc_sdram_inti_p1_ras_n <= 1'd1;
	videosoc_sdram_inti_p1_we_n <= 1'd1;
	if (videosoc_sdram_phaseinjector1_command_issue_re) begin
		videosoc_sdram_inti_p1_cs_n <= (~videosoc_sdram_phaseinjector1_command_storage[0]);
		videosoc_sdram_inti_p1_we_n <= (~videosoc_sdram_phaseinjector1_command_storage[1]);
		videosoc_sdram_inti_p1_cas_n <= (~videosoc_sdram_phaseinjector1_command_storage[2]);
		videosoc_sdram_inti_p1_ras_n <= (~videosoc_sdram_phaseinjector1_command_storage[3]);
	end else begin
		videosoc_sdram_inti_p1_cs_n <= 1'd1;
		videosoc_sdram_inti_p1_we_n <= 1'd1;
		videosoc_sdram_inti_p1_cas_n <= 1'd1;
		videosoc_sdram_inti_p1_ras_n <= 1'd1;
	end
end
assign videosoc_sdram_inti_p1_address = videosoc_sdram_phaseinjector1_address_storage;
assign videosoc_sdram_inti_p1_bank = videosoc_sdram_phaseinjector1_baddress_storage;
assign videosoc_sdram_inti_p1_wrdata_en = (videosoc_sdram_phaseinjector1_command_issue_re & videosoc_sdram_phaseinjector1_command_storage[4]);
assign videosoc_sdram_inti_p1_rddata_en = (videosoc_sdram_phaseinjector1_command_issue_re & videosoc_sdram_phaseinjector1_command_storage[5]);
assign videosoc_sdram_inti_p1_wrdata = videosoc_sdram_phaseinjector1_wrdata_storage;
assign videosoc_sdram_inti_p1_wrdata_mask = 1'd0;
always @(*) begin
	videosoc_sdram_inti_p2_cs_n <= 1'd1;
	videosoc_sdram_inti_p2_ras_n <= 1'd1;
	videosoc_sdram_inti_p2_we_n <= 1'd1;
	videosoc_sdram_inti_p2_cas_n <= 1'd1;
	if (videosoc_sdram_phaseinjector2_command_issue_re) begin
		videosoc_sdram_inti_p2_cs_n <= (~videosoc_sdram_phaseinjector2_command_storage[0]);
		videosoc_sdram_inti_p2_we_n <= (~videosoc_sdram_phaseinjector2_command_storage[1]);
		videosoc_sdram_inti_p2_cas_n <= (~videosoc_sdram_phaseinjector2_command_storage[2]);
		videosoc_sdram_inti_p2_ras_n <= (~videosoc_sdram_phaseinjector2_command_storage[3]);
	end else begin
		videosoc_sdram_inti_p2_cs_n <= 1'd1;
		videosoc_sdram_inti_p2_we_n <= 1'd1;
		videosoc_sdram_inti_p2_cas_n <= 1'd1;
		videosoc_sdram_inti_p2_ras_n <= 1'd1;
	end
end
assign videosoc_sdram_inti_p2_address = videosoc_sdram_phaseinjector2_address_storage;
assign videosoc_sdram_inti_p2_bank = videosoc_sdram_phaseinjector2_baddress_storage;
assign videosoc_sdram_inti_p2_wrdata_en = (videosoc_sdram_phaseinjector2_command_issue_re & videosoc_sdram_phaseinjector2_command_storage[4]);
assign videosoc_sdram_inti_p2_rddata_en = (videosoc_sdram_phaseinjector2_command_issue_re & videosoc_sdram_phaseinjector2_command_storage[5]);
assign videosoc_sdram_inti_p2_wrdata = videosoc_sdram_phaseinjector2_wrdata_storage;
assign videosoc_sdram_inti_p2_wrdata_mask = 1'd0;
always @(*) begin
	videosoc_sdram_inti_p3_ras_n <= 1'd1;
	videosoc_sdram_inti_p3_we_n <= 1'd1;
	videosoc_sdram_inti_p3_cas_n <= 1'd1;
	videosoc_sdram_inti_p3_cs_n <= 1'd1;
	if (videosoc_sdram_phaseinjector3_command_issue_re) begin
		videosoc_sdram_inti_p3_cs_n <= (~videosoc_sdram_phaseinjector3_command_storage[0]);
		videosoc_sdram_inti_p3_we_n <= (~videosoc_sdram_phaseinjector3_command_storage[1]);
		videosoc_sdram_inti_p3_cas_n <= (~videosoc_sdram_phaseinjector3_command_storage[2]);
		videosoc_sdram_inti_p3_ras_n <= (~videosoc_sdram_phaseinjector3_command_storage[3]);
	end else begin
		videosoc_sdram_inti_p3_cs_n <= 1'd1;
		videosoc_sdram_inti_p3_we_n <= 1'd1;
		videosoc_sdram_inti_p3_cas_n <= 1'd1;
		videosoc_sdram_inti_p3_ras_n <= 1'd1;
	end
end
assign videosoc_sdram_inti_p3_address = videosoc_sdram_phaseinjector3_address_storage;
assign videosoc_sdram_inti_p3_bank = videosoc_sdram_phaseinjector3_baddress_storage;
assign videosoc_sdram_inti_p3_wrdata_en = (videosoc_sdram_phaseinjector3_command_issue_re & videosoc_sdram_phaseinjector3_command_storage[4]);
assign videosoc_sdram_inti_p3_rddata_en = (videosoc_sdram_phaseinjector3_command_issue_re & videosoc_sdram_phaseinjector3_command_storage[5]);
assign videosoc_sdram_inti_p3_wrdata = videosoc_sdram_phaseinjector3_wrdata_storage;
assign videosoc_sdram_inti_p3_wrdata_mask = 1'd0;
assign videosoc_sdram_bankmachine0_req_valid = videosoc_sdram_interface_bank0_valid;
assign videosoc_sdram_interface_bank0_ready = videosoc_sdram_bankmachine0_req_ready;
assign videosoc_sdram_bankmachine0_req_we = videosoc_sdram_interface_bank0_we;
assign videosoc_sdram_bankmachine0_req_adr = videosoc_sdram_interface_bank0_adr;
assign videosoc_sdram_interface_bank0_lock = videosoc_sdram_bankmachine0_req_lock;
assign videosoc_sdram_interface_bank0_wdata_ready = videosoc_sdram_bankmachine0_req_wdata_ready;
assign videosoc_sdram_interface_bank0_rdata_valid = videosoc_sdram_bankmachine0_req_rdata_valid;
assign videosoc_sdram_bankmachine1_req_valid = videosoc_sdram_interface_bank1_valid;
assign videosoc_sdram_interface_bank1_ready = videosoc_sdram_bankmachine1_req_ready;
assign videosoc_sdram_bankmachine1_req_we = videosoc_sdram_interface_bank1_we;
assign videosoc_sdram_bankmachine1_req_adr = videosoc_sdram_interface_bank1_adr;
assign videosoc_sdram_interface_bank1_lock = videosoc_sdram_bankmachine1_req_lock;
assign videosoc_sdram_interface_bank1_wdata_ready = videosoc_sdram_bankmachine1_req_wdata_ready;
assign videosoc_sdram_interface_bank1_rdata_valid = videosoc_sdram_bankmachine1_req_rdata_valid;
assign videosoc_sdram_bankmachine2_req_valid = videosoc_sdram_interface_bank2_valid;
assign videosoc_sdram_interface_bank2_ready = videosoc_sdram_bankmachine2_req_ready;
assign videosoc_sdram_bankmachine2_req_we = videosoc_sdram_interface_bank2_we;
assign videosoc_sdram_bankmachine2_req_adr = videosoc_sdram_interface_bank2_adr;
assign videosoc_sdram_interface_bank2_lock = videosoc_sdram_bankmachine2_req_lock;
assign videosoc_sdram_interface_bank2_wdata_ready = videosoc_sdram_bankmachine2_req_wdata_ready;
assign videosoc_sdram_interface_bank2_rdata_valid = videosoc_sdram_bankmachine2_req_rdata_valid;
assign videosoc_sdram_bankmachine3_req_valid = videosoc_sdram_interface_bank3_valid;
assign videosoc_sdram_interface_bank3_ready = videosoc_sdram_bankmachine3_req_ready;
assign videosoc_sdram_bankmachine3_req_we = videosoc_sdram_interface_bank3_we;
assign videosoc_sdram_bankmachine3_req_adr = videosoc_sdram_interface_bank3_adr;
assign videosoc_sdram_interface_bank3_lock = videosoc_sdram_bankmachine3_req_lock;
assign videosoc_sdram_interface_bank3_wdata_ready = videosoc_sdram_bankmachine3_req_wdata_ready;
assign videosoc_sdram_interface_bank3_rdata_valid = videosoc_sdram_bankmachine3_req_rdata_valid;
assign videosoc_sdram_bankmachine4_req_valid = videosoc_sdram_interface_bank4_valid;
assign videosoc_sdram_interface_bank4_ready = videosoc_sdram_bankmachine4_req_ready;
assign videosoc_sdram_bankmachine4_req_we = videosoc_sdram_interface_bank4_we;
assign videosoc_sdram_bankmachine4_req_adr = videosoc_sdram_interface_bank4_adr;
assign videosoc_sdram_interface_bank4_lock = videosoc_sdram_bankmachine4_req_lock;
assign videosoc_sdram_interface_bank4_wdata_ready = videosoc_sdram_bankmachine4_req_wdata_ready;
assign videosoc_sdram_interface_bank4_rdata_valid = videosoc_sdram_bankmachine4_req_rdata_valid;
assign videosoc_sdram_bankmachine5_req_valid = videosoc_sdram_interface_bank5_valid;
assign videosoc_sdram_interface_bank5_ready = videosoc_sdram_bankmachine5_req_ready;
assign videosoc_sdram_bankmachine5_req_we = videosoc_sdram_interface_bank5_we;
assign videosoc_sdram_bankmachine5_req_adr = videosoc_sdram_interface_bank5_adr;
assign videosoc_sdram_interface_bank5_lock = videosoc_sdram_bankmachine5_req_lock;
assign videosoc_sdram_interface_bank5_wdata_ready = videosoc_sdram_bankmachine5_req_wdata_ready;
assign videosoc_sdram_interface_bank5_rdata_valid = videosoc_sdram_bankmachine5_req_rdata_valid;
assign videosoc_sdram_bankmachine6_req_valid = videosoc_sdram_interface_bank6_valid;
assign videosoc_sdram_interface_bank6_ready = videosoc_sdram_bankmachine6_req_ready;
assign videosoc_sdram_bankmachine6_req_we = videosoc_sdram_interface_bank6_we;
assign videosoc_sdram_bankmachine6_req_adr = videosoc_sdram_interface_bank6_adr;
assign videosoc_sdram_interface_bank6_lock = videosoc_sdram_bankmachine6_req_lock;
assign videosoc_sdram_interface_bank6_wdata_ready = videosoc_sdram_bankmachine6_req_wdata_ready;
assign videosoc_sdram_interface_bank6_rdata_valid = videosoc_sdram_bankmachine6_req_rdata_valid;
assign videosoc_sdram_bankmachine7_req_valid = videosoc_sdram_interface_bank7_valid;
assign videosoc_sdram_interface_bank7_ready = videosoc_sdram_bankmachine7_req_ready;
assign videosoc_sdram_bankmachine7_req_we = videosoc_sdram_interface_bank7_we;
assign videosoc_sdram_bankmachine7_req_adr = videosoc_sdram_interface_bank7_adr;
assign videosoc_sdram_interface_bank7_lock = videosoc_sdram_bankmachine7_req_lock;
assign videosoc_sdram_interface_bank7_wdata_ready = videosoc_sdram_bankmachine7_req_wdata_ready;
assign videosoc_sdram_interface_bank7_rdata_valid = videosoc_sdram_bankmachine7_req_rdata_valid;
assign videosoc_sdram_wait = (1'd1 & (~videosoc_sdram_done));
assign videosoc_sdram_done = (videosoc_sdram_count == 1'd0);
always @(*) begin
	videosoc_sdram_seq_start <= 1'd0;
	refresher_next_state <= 2'd0;
	videosoc_sdram_cmd_last <= 1'd0;
	videosoc_sdram_cmd_valid <= 1'd0;
	refresher_next_state <= refresher_state;
	case (refresher_state)
		1'd1: begin
			videosoc_sdram_cmd_valid <= 1'd1;
			if (videosoc_sdram_cmd_ready) begin
				videosoc_sdram_seq_start <= 1'd1;
				refresher_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (videosoc_sdram_seq_done) begin
				videosoc_sdram_cmd_last <= 1'd1;
				refresher_next_state <= 1'd0;
			end else begin
				videosoc_sdram_cmd_valid <= 1'd1;
			end
		end
		default: begin
			if (videosoc_sdram_done) begin
				refresher_next_state <= 1'd1;
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine0_sink_valid = videosoc_sdram_bankmachine0_req_valid;
assign videosoc_sdram_bankmachine0_req_ready = videosoc_sdram_bankmachine0_sink_ready;
assign videosoc_sdram_bankmachine0_sink_payload_we = videosoc_sdram_bankmachine0_req_we;
assign videosoc_sdram_bankmachine0_sink_payload_adr = videosoc_sdram_bankmachine0_req_adr;
assign videosoc_sdram_bankmachine0_source_ready = (videosoc_sdram_bankmachine0_req_wdata_ready | videosoc_sdram_bankmachine0_req_rdata_valid);
assign videosoc_sdram_bankmachine0_req_lock = videosoc_sdram_bankmachine0_source_valid;
assign videosoc_sdram_bankmachine0_hit = (videosoc_sdram_bankmachine0_openrow == videosoc_sdram_bankmachine0_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine0_cmd_payload_ba = 1'd0;
always @(*) begin
	videosoc_sdram_bankmachine0_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine0_sel_row_adr) begin
		videosoc_sdram_bankmachine0_cmd_payload_a <= videosoc_sdram_bankmachine0_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine0_cmd_payload_a <= {videosoc_sdram_bankmachine0_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine0_wait = (~((videosoc_sdram_bankmachine0_cmd_valid & videosoc_sdram_bankmachine0_cmd_ready) & videosoc_sdram_bankmachine0_cmd_payload_is_write));
assign videosoc_sdram_bankmachine0_syncfifo0_din = {videosoc_sdram_bankmachine0_fifo_in_last, videosoc_sdram_bankmachine0_fifo_in_first, videosoc_sdram_bankmachine0_fifo_in_payload_adr, videosoc_sdram_bankmachine0_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine0_fifo_out_last, videosoc_sdram_bankmachine0_fifo_out_first, videosoc_sdram_bankmachine0_fifo_out_payload_adr, videosoc_sdram_bankmachine0_fifo_out_payload_we} = videosoc_sdram_bankmachine0_syncfifo0_dout;
assign videosoc_sdram_bankmachine0_sink_ready = videosoc_sdram_bankmachine0_syncfifo0_writable;
assign videosoc_sdram_bankmachine0_syncfifo0_we = videosoc_sdram_bankmachine0_sink_valid;
assign videosoc_sdram_bankmachine0_fifo_in_first = videosoc_sdram_bankmachine0_sink_first;
assign videosoc_sdram_bankmachine0_fifo_in_last = videosoc_sdram_bankmachine0_sink_last;
assign videosoc_sdram_bankmachine0_fifo_in_payload_we = videosoc_sdram_bankmachine0_sink_payload_we;
assign videosoc_sdram_bankmachine0_fifo_in_payload_adr = videosoc_sdram_bankmachine0_sink_payload_adr;
assign videosoc_sdram_bankmachine0_source_valid = videosoc_sdram_bankmachine0_syncfifo0_readable;
assign videosoc_sdram_bankmachine0_source_first = videosoc_sdram_bankmachine0_fifo_out_first;
assign videosoc_sdram_bankmachine0_source_last = videosoc_sdram_bankmachine0_fifo_out_last;
assign videosoc_sdram_bankmachine0_source_payload_we = videosoc_sdram_bankmachine0_fifo_out_payload_we;
assign videosoc_sdram_bankmachine0_source_payload_adr = videosoc_sdram_bankmachine0_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine0_syncfifo0_re = videosoc_sdram_bankmachine0_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine0_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine0_replace) begin
		videosoc_sdram_bankmachine0_wrport_adr <= (videosoc_sdram_bankmachine0_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine0_wrport_adr <= videosoc_sdram_bankmachine0_produce;
	end
end
assign videosoc_sdram_bankmachine0_wrport_dat_w = videosoc_sdram_bankmachine0_syncfifo0_din;
assign videosoc_sdram_bankmachine0_wrport_we = (videosoc_sdram_bankmachine0_syncfifo0_we & (videosoc_sdram_bankmachine0_syncfifo0_writable | videosoc_sdram_bankmachine0_replace));
assign videosoc_sdram_bankmachine0_do_read = (videosoc_sdram_bankmachine0_syncfifo0_readable & videosoc_sdram_bankmachine0_syncfifo0_re);
assign videosoc_sdram_bankmachine0_rdport_adr = videosoc_sdram_bankmachine0_consume;
assign videosoc_sdram_bankmachine0_syncfifo0_dout = videosoc_sdram_bankmachine0_rdport_dat_r;
assign videosoc_sdram_bankmachine0_syncfifo0_writable = (videosoc_sdram_bankmachine0_level != 4'd8);
assign videosoc_sdram_bankmachine0_syncfifo0_readable = (videosoc_sdram_bankmachine0_level != 1'd0);
assign videosoc_sdram_bankmachine0_done = (videosoc_sdram_bankmachine0_count == 1'd0);
always @(*) begin
	videosoc_sdram_bankmachine0_track_open <= 1'd0;
	videosoc_sdram_bankmachine0_track_close <= 1'd0;
	videosoc_sdram_bankmachine0_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine0_cmd_payload_ras <= 1'd0;
	videosoc_sdram_bankmachine0_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine0_sel_row_adr <= 1'd0;
	videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd0;
	videosoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine0_req_wdata_ready <= 1'd0;
	videosoc_sdram_bankmachine0_req_rdata_valid <= 1'd0;
	videosoc_sdram_bankmachine0_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine0_cmd_valid <= 1'd0;
	bankmachine0_next_state <= 3'd0;
	bankmachine0_next_state <= bankmachine0_state;
	case (bankmachine0_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine0_done) begin
				videosoc_sdram_bankmachine0_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine0_cmd_ready) begin
					bankmachine0_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine0_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine0_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine0_track_open <= 1'd1;
			videosoc_sdram_bankmachine0_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine0_cmd_ready) begin
				bankmachine0_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine0_done) begin
				videosoc_sdram_bankmachine0_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine0_track_close <= 1'd1;
			videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine0_refresh_req)) begin
				bankmachine0_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine0_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine0_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine0_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine0_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine0_refresh_req) begin
				bankmachine0_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine0_source_valid) begin
					if (videosoc_sdram_bankmachine0_has_openrow) begin
						if (videosoc_sdram_bankmachine0_hit) begin
							videosoc_sdram_bankmachine0_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine0_source_payload_we) begin
								videosoc_sdram_bankmachine0_req_wdata_ready <= videosoc_sdram_bankmachine0_cmd_ready;
								videosoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine0_req_rdata_valid <= videosoc_sdram_bankmachine0_cmd_ready;
								videosoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine0_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine0_next_state <= 1'd1;
						end
					end else begin
						bankmachine0_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine1_sink_valid = videosoc_sdram_bankmachine1_req_valid;
assign videosoc_sdram_bankmachine1_req_ready = videosoc_sdram_bankmachine1_sink_ready;
assign videosoc_sdram_bankmachine1_sink_payload_we = videosoc_sdram_bankmachine1_req_we;
assign videosoc_sdram_bankmachine1_sink_payload_adr = videosoc_sdram_bankmachine1_req_adr;
assign videosoc_sdram_bankmachine1_source_ready = (videosoc_sdram_bankmachine1_req_wdata_ready | videosoc_sdram_bankmachine1_req_rdata_valid);
assign videosoc_sdram_bankmachine1_req_lock = videosoc_sdram_bankmachine1_source_valid;
assign videosoc_sdram_bankmachine1_hit = (videosoc_sdram_bankmachine1_openrow == videosoc_sdram_bankmachine1_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine1_cmd_payload_ba = 1'd1;
always @(*) begin
	videosoc_sdram_bankmachine1_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine1_sel_row_adr) begin
		videosoc_sdram_bankmachine1_cmd_payload_a <= videosoc_sdram_bankmachine1_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine1_cmd_payload_a <= {videosoc_sdram_bankmachine1_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine1_wait = (~((videosoc_sdram_bankmachine1_cmd_valid & videosoc_sdram_bankmachine1_cmd_ready) & videosoc_sdram_bankmachine1_cmd_payload_is_write));
assign videosoc_sdram_bankmachine1_syncfifo1_din = {videosoc_sdram_bankmachine1_fifo_in_last, videosoc_sdram_bankmachine1_fifo_in_first, videosoc_sdram_bankmachine1_fifo_in_payload_adr, videosoc_sdram_bankmachine1_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine1_fifo_out_last, videosoc_sdram_bankmachine1_fifo_out_first, videosoc_sdram_bankmachine1_fifo_out_payload_adr, videosoc_sdram_bankmachine1_fifo_out_payload_we} = videosoc_sdram_bankmachine1_syncfifo1_dout;
assign videosoc_sdram_bankmachine1_sink_ready = videosoc_sdram_bankmachine1_syncfifo1_writable;
assign videosoc_sdram_bankmachine1_syncfifo1_we = videosoc_sdram_bankmachine1_sink_valid;
assign videosoc_sdram_bankmachine1_fifo_in_first = videosoc_sdram_bankmachine1_sink_first;
assign videosoc_sdram_bankmachine1_fifo_in_last = videosoc_sdram_bankmachine1_sink_last;
assign videosoc_sdram_bankmachine1_fifo_in_payload_we = videosoc_sdram_bankmachine1_sink_payload_we;
assign videosoc_sdram_bankmachine1_fifo_in_payload_adr = videosoc_sdram_bankmachine1_sink_payload_adr;
assign videosoc_sdram_bankmachine1_source_valid = videosoc_sdram_bankmachine1_syncfifo1_readable;
assign videosoc_sdram_bankmachine1_source_first = videosoc_sdram_bankmachine1_fifo_out_first;
assign videosoc_sdram_bankmachine1_source_last = videosoc_sdram_bankmachine1_fifo_out_last;
assign videosoc_sdram_bankmachine1_source_payload_we = videosoc_sdram_bankmachine1_fifo_out_payload_we;
assign videosoc_sdram_bankmachine1_source_payload_adr = videosoc_sdram_bankmachine1_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine1_syncfifo1_re = videosoc_sdram_bankmachine1_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine1_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine1_replace) begin
		videosoc_sdram_bankmachine1_wrport_adr <= (videosoc_sdram_bankmachine1_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine1_wrport_adr <= videosoc_sdram_bankmachine1_produce;
	end
end
assign videosoc_sdram_bankmachine1_wrport_dat_w = videosoc_sdram_bankmachine1_syncfifo1_din;
assign videosoc_sdram_bankmachine1_wrport_we = (videosoc_sdram_bankmachine1_syncfifo1_we & (videosoc_sdram_bankmachine1_syncfifo1_writable | videosoc_sdram_bankmachine1_replace));
assign videosoc_sdram_bankmachine1_do_read = (videosoc_sdram_bankmachine1_syncfifo1_readable & videosoc_sdram_bankmachine1_syncfifo1_re);
assign videosoc_sdram_bankmachine1_rdport_adr = videosoc_sdram_bankmachine1_consume;
assign videosoc_sdram_bankmachine1_syncfifo1_dout = videosoc_sdram_bankmachine1_rdport_dat_r;
assign videosoc_sdram_bankmachine1_syncfifo1_writable = (videosoc_sdram_bankmachine1_level != 4'd8);
assign videosoc_sdram_bankmachine1_syncfifo1_readable = (videosoc_sdram_bankmachine1_level != 1'd0);
assign videosoc_sdram_bankmachine1_done = (videosoc_sdram_bankmachine1_count == 1'd0);
always @(*) begin
	videosoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine1_req_wdata_ready <= 1'd0;
	videosoc_sdram_bankmachine1_req_rdata_valid <= 1'd0;
	videosoc_sdram_bankmachine1_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine1_cmd_valid <= 1'd0;
	videosoc_sdram_bankmachine1_track_open <= 1'd0;
	videosoc_sdram_bankmachine1_track_close <= 1'd0;
	videosoc_sdram_bankmachine1_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine1_cmd_payload_ras <= 1'd0;
	bankmachine1_next_state <= 3'd0;
	videosoc_sdram_bankmachine1_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine1_sel_row_adr <= 1'd0;
	videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd0;
	bankmachine1_next_state <= bankmachine1_state;
	case (bankmachine1_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine1_done) begin
				videosoc_sdram_bankmachine1_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine1_cmd_ready) begin
					bankmachine1_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine1_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine1_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine1_track_open <= 1'd1;
			videosoc_sdram_bankmachine1_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine1_cmd_ready) begin
				bankmachine1_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine1_done) begin
				videosoc_sdram_bankmachine1_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine1_track_close <= 1'd1;
			videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine1_refresh_req)) begin
				bankmachine1_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine1_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine1_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine1_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine1_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine1_refresh_req) begin
				bankmachine1_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine1_source_valid) begin
					if (videosoc_sdram_bankmachine1_has_openrow) begin
						if (videosoc_sdram_bankmachine1_hit) begin
							videosoc_sdram_bankmachine1_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine1_source_payload_we) begin
								videosoc_sdram_bankmachine1_req_wdata_ready <= videosoc_sdram_bankmachine1_cmd_ready;
								videosoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine1_req_rdata_valid <= videosoc_sdram_bankmachine1_cmd_ready;
								videosoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine1_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine1_next_state <= 1'd1;
						end
					end else begin
						bankmachine1_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine2_sink_valid = videosoc_sdram_bankmachine2_req_valid;
assign videosoc_sdram_bankmachine2_req_ready = videosoc_sdram_bankmachine2_sink_ready;
assign videosoc_sdram_bankmachine2_sink_payload_we = videosoc_sdram_bankmachine2_req_we;
assign videosoc_sdram_bankmachine2_sink_payload_adr = videosoc_sdram_bankmachine2_req_adr;
assign videosoc_sdram_bankmachine2_source_ready = (videosoc_sdram_bankmachine2_req_wdata_ready | videosoc_sdram_bankmachine2_req_rdata_valid);
assign videosoc_sdram_bankmachine2_req_lock = videosoc_sdram_bankmachine2_source_valid;
assign videosoc_sdram_bankmachine2_hit = (videosoc_sdram_bankmachine2_openrow == videosoc_sdram_bankmachine2_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine2_cmd_payload_ba = 2'd2;
always @(*) begin
	videosoc_sdram_bankmachine2_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine2_sel_row_adr) begin
		videosoc_sdram_bankmachine2_cmd_payload_a <= videosoc_sdram_bankmachine2_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine2_cmd_payload_a <= {videosoc_sdram_bankmachine2_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine2_wait = (~((videosoc_sdram_bankmachine2_cmd_valid & videosoc_sdram_bankmachine2_cmd_ready) & videosoc_sdram_bankmachine2_cmd_payload_is_write));
assign videosoc_sdram_bankmachine2_syncfifo2_din = {videosoc_sdram_bankmachine2_fifo_in_last, videosoc_sdram_bankmachine2_fifo_in_first, videosoc_sdram_bankmachine2_fifo_in_payload_adr, videosoc_sdram_bankmachine2_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine2_fifo_out_last, videosoc_sdram_bankmachine2_fifo_out_first, videosoc_sdram_bankmachine2_fifo_out_payload_adr, videosoc_sdram_bankmachine2_fifo_out_payload_we} = videosoc_sdram_bankmachine2_syncfifo2_dout;
assign videosoc_sdram_bankmachine2_sink_ready = videosoc_sdram_bankmachine2_syncfifo2_writable;
assign videosoc_sdram_bankmachine2_syncfifo2_we = videosoc_sdram_bankmachine2_sink_valid;
assign videosoc_sdram_bankmachine2_fifo_in_first = videosoc_sdram_bankmachine2_sink_first;
assign videosoc_sdram_bankmachine2_fifo_in_last = videosoc_sdram_bankmachine2_sink_last;
assign videosoc_sdram_bankmachine2_fifo_in_payload_we = videosoc_sdram_bankmachine2_sink_payload_we;
assign videosoc_sdram_bankmachine2_fifo_in_payload_adr = videosoc_sdram_bankmachine2_sink_payload_adr;
assign videosoc_sdram_bankmachine2_source_valid = videosoc_sdram_bankmachine2_syncfifo2_readable;
assign videosoc_sdram_bankmachine2_source_first = videosoc_sdram_bankmachine2_fifo_out_first;
assign videosoc_sdram_bankmachine2_source_last = videosoc_sdram_bankmachine2_fifo_out_last;
assign videosoc_sdram_bankmachine2_source_payload_we = videosoc_sdram_bankmachine2_fifo_out_payload_we;
assign videosoc_sdram_bankmachine2_source_payload_adr = videosoc_sdram_bankmachine2_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine2_syncfifo2_re = videosoc_sdram_bankmachine2_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine2_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine2_replace) begin
		videosoc_sdram_bankmachine2_wrport_adr <= (videosoc_sdram_bankmachine2_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine2_wrport_adr <= videosoc_sdram_bankmachine2_produce;
	end
end
assign videosoc_sdram_bankmachine2_wrport_dat_w = videosoc_sdram_bankmachine2_syncfifo2_din;
assign videosoc_sdram_bankmachine2_wrport_we = (videosoc_sdram_bankmachine2_syncfifo2_we & (videosoc_sdram_bankmachine2_syncfifo2_writable | videosoc_sdram_bankmachine2_replace));
assign videosoc_sdram_bankmachine2_do_read = (videosoc_sdram_bankmachine2_syncfifo2_readable & videosoc_sdram_bankmachine2_syncfifo2_re);
assign videosoc_sdram_bankmachine2_rdport_adr = videosoc_sdram_bankmachine2_consume;
assign videosoc_sdram_bankmachine2_syncfifo2_dout = videosoc_sdram_bankmachine2_rdport_dat_r;
assign videosoc_sdram_bankmachine2_syncfifo2_writable = (videosoc_sdram_bankmachine2_level != 4'd8);
assign videosoc_sdram_bankmachine2_syncfifo2_readable = (videosoc_sdram_bankmachine2_level != 1'd0);
assign videosoc_sdram_bankmachine2_done = (videosoc_sdram_bankmachine2_count == 1'd0);
always @(*) begin
	videosoc_sdram_bankmachine2_track_open <= 1'd0;
	videosoc_sdram_bankmachine2_track_close <= 1'd0;
	videosoc_sdram_bankmachine2_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine2_cmd_payload_ras <= 1'd0;
	videosoc_sdram_bankmachine2_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine2_sel_row_adr <= 1'd0;
	videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd0;
	videosoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine2_req_wdata_ready <= 1'd0;
	videosoc_sdram_bankmachine2_req_rdata_valid <= 1'd0;
	bankmachine2_next_state <= 3'd0;
	videosoc_sdram_bankmachine2_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine2_cmd_valid <= 1'd0;
	bankmachine2_next_state <= bankmachine2_state;
	case (bankmachine2_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine2_done) begin
				videosoc_sdram_bankmachine2_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine2_cmd_ready) begin
					bankmachine2_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine2_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine2_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine2_track_open <= 1'd1;
			videosoc_sdram_bankmachine2_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine2_cmd_ready) begin
				bankmachine2_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine2_done) begin
				videosoc_sdram_bankmachine2_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine2_track_close <= 1'd1;
			videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine2_refresh_req)) begin
				bankmachine2_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine2_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine2_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine2_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine2_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine2_refresh_req) begin
				bankmachine2_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine2_source_valid) begin
					if (videosoc_sdram_bankmachine2_has_openrow) begin
						if (videosoc_sdram_bankmachine2_hit) begin
							videosoc_sdram_bankmachine2_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine2_source_payload_we) begin
								videosoc_sdram_bankmachine2_req_wdata_ready <= videosoc_sdram_bankmachine2_cmd_ready;
								videosoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine2_req_rdata_valid <= videosoc_sdram_bankmachine2_cmd_ready;
								videosoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine2_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine2_next_state <= 1'd1;
						end
					end else begin
						bankmachine2_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine3_sink_valid = videosoc_sdram_bankmachine3_req_valid;
assign videosoc_sdram_bankmachine3_req_ready = videosoc_sdram_bankmachine3_sink_ready;
assign videosoc_sdram_bankmachine3_sink_payload_we = videosoc_sdram_bankmachine3_req_we;
assign videosoc_sdram_bankmachine3_sink_payload_adr = videosoc_sdram_bankmachine3_req_adr;
assign videosoc_sdram_bankmachine3_source_ready = (videosoc_sdram_bankmachine3_req_wdata_ready | videosoc_sdram_bankmachine3_req_rdata_valid);
assign videosoc_sdram_bankmachine3_req_lock = videosoc_sdram_bankmachine3_source_valid;
assign videosoc_sdram_bankmachine3_hit = (videosoc_sdram_bankmachine3_openrow == videosoc_sdram_bankmachine3_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine3_cmd_payload_ba = 2'd3;
always @(*) begin
	videosoc_sdram_bankmachine3_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine3_sel_row_adr) begin
		videosoc_sdram_bankmachine3_cmd_payload_a <= videosoc_sdram_bankmachine3_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine3_cmd_payload_a <= {videosoc_sdram_bankmachine3_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine3_wait = (~((videosoc_sdram_bankmachine3_cmd_valid & videosoc_sdram_bankmachine3_cmd_ready) & videosoc_sdram_bankmachine3_cmd_payload_is_write));
assign videosoc_sdram_bankmachine3_syncfifo3_din = {videosoc_sdram_bankmachine3_fifo_in_last, videosoc_sdram_bankmachine3_fifo_in_first, videosoc_sdram_bankmachine3_fifo_in_payload_adr, videosoc_sdram_bankmachine3_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine3_fifo_out_last, videosoc_sdram_bankmachine3_fifo_out_first, videosoc_sdram_bankmachine3_fifo_out_payload_adr, videosoc_sdram_bankmachine3_fifo_out_payload_we} = videosoc_sdram_bankmachine3_syncfifo3_dout;
assign videosoc_sdram_bankmachine3_sink_ready = videosoc_sdram_bankmachine3_syncfifo3_writable;
assign videosoc_sdram_bankmachine3_syncfifo3_we = videosoc_sdram_bankmachine3_sink_valid;
assign videosoc_sdram_bankmachine3_fifo_in_first = videosoc_sdram_bankmachine3_sink_first;
assign videosoc_sdram_bankmachine3_fifo_in_last = videosoc_sdram_bankmachine3_sink_last;
assign videosoc_sdram_bankmachine3_fifo_in_payload_we = videosoc_sdram_bankmachine3_sink_payload_we;
assign videosoc_sdram_bankmachine3_fifo_in_payload_adr = videosoc_sdram_bankmachine3_sink_payload_adr;
assign videosoc_sdram_bankmachine3_source_valid = videosoc_sdram_bankmachine3_syncfifo3_readable;
assign videosoc_sdram_bankmachine3_source_first = videosoc_sdram_bankmachine3_fifo_out_first;
assign videosoc_sdram_bankmachine3_source_last = videosoc_sdram_bankmachine3_fifo_out_last;
assign videosoc_sdram_bankmachine3_source_payload_we = videosoc_sdram_bankmachine3_fifo_out_payload_we;
assign videosoc_sdram_bankmachine3_source_payload_adr = videosoc_sdram_bankmachine3_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine3_syncfifo3_re = videosoc_sdram_bankmachine3_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine3_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine3_replace) begin
		videosoc_sdram_bankmachine3_wrport_adr <= (videosoc_sdram_bankmachine3_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine3_wrport_adr <= videosoc_sdram_bankmachine3_produce;
	end
end
assign videosoc_sdram_bankmachine3_wrport_dat_w = videosoc_sdram_bankmachine3_syncfifo3_din;
assign videosoc_sdram_bankmachine3_wrport_we = (videosoc_sdram_bankmachine3_syncfifo3_we & (videosoc_sdram_bankmachine3_syncfifo3_writable | videosoc_sdram_bankmachine3_replace));
assign videosoc_sdram_bankmachine3_do_read = (videosoc_sdram_bankmachine3_syncfifo3_readable & videosoc_sdram_bankmachine3_syncfifo3_re);
assign videosoc_sdram_bankmachine3_rdport_adr = videosoc_sdram_bankmachine3_consume;
assign videosoc_sdram_bankmachine3_syncfifo3_dout = videosoc_sdram_bankmachine3_rdport_dat_r;
assign videosoc_sdram_bankmachine3_syncfifo3_writable = (videosoc_sdram_bankmachine3_level != 4'd8);
assign videosoc_sdram_bankmachine3_syncfifo3_readable = (videosoc_sdram_bankmachine3_level != 1'd0);
assign videosoc_sdram_bankmachine3_done = (videosoc_sdram_bankmachine3_count == 1'd0);
always @(*) begin
	videosoc_sdram_bankmachine3_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine3_cmd_valid <= 1'd0;
	videosoc_sdram_bankmachine3_track_open <= 1'd0;
	bankmachine3_next_state <= 3'd0;
	videosoc_sdram_bankmachine3_track_close <= 1'd0;
	videosoc_sdram_bankmachine3_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine3_cmd_payload_ras <= 1'd0;
	videosoc_sdram_bankmachine3_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine3_sel_row_adr <= 1'd0;
	videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd0;
	videosoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine3_req_wdata_ready <= 1'd0;
	videosoc_sdram_bankmachine3_req_rdata_valid <= 1'd0;
	bankmachine3_next_state <= bankmachine3_state;
	case (bankmachine3_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine3_done) begin
				videosoc_sdram_bankmachine3_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine3_cmd_ready) begin
					bankmachine3_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine3_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine3_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine3_track_open <= 1'd1;
			videosoc_sdram_bankmachine3_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine3_cmd_ready) begin
				bankmachine3_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine3_done) begin
				videosoc_sdram_bankmachine3_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine3_track_close <= 1'd1;
			videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine3_refresh_req)) begin
				bankmachine3_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine3_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine3_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine3_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine3_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine3_refresh_req) begin
				bankmachine3_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine3_source_valid) begin
					if (videosoc_sdram_bankmachine3_has_openrow) begin
						if (videosoc_sdram_bankmachine3_hit) begin
							videosoc_sdram_bankmachine3_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine3_source_payload_we) begin
								videosoc_sdram_bankmachine3_req_wdata_ready <= videosoc_sdram_bankmachine3_cmd_ready;
								videosoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine3_req_rdata_valid <= videosoc_sdram_bankmachine3_cmd_ready;
								videosoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine3_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine3_next_state <= 1'd1;
						end
					end else begin
						bankmachine3_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine4_sink_valid = videosoc_sdram_bankmachine4_req_valid;
assign videosoc_sdram_bankmachine4_req_ready = videosoc_sdram_bankmachine4_sink_ready;
assign videosoc_sdram_bankmachine4_sink_payload_we = videosoc_sdram_bankmachine4_req_we;
assign videosoc_sdram_bankmachine4_sink_payload_adr = videosoc_sdram_bankmachine4_req_adr;
assign videosoc_sdram_bankmachine4_source_ready = (videosoc_sdram_bankmachine4_req_wdata_ready | videosoc_sdram_bankmachine4_req_rdata_valid);
assign videosoc_sdram_bankmachine4_req_lock = videosoc_sdram_bankmachine4_source_valid;
assign videosoc_sdram_bankmachine4_hit = (videosoc_sdram_bankmachine4_openrow == videosoc_sdram_bankmachine4_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine4_cmd_payload_ba = 3'd4;
always @(*) begin
	videosoc_sdram_bankmachine4_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine4_sel_row_adr) begin
		videosoc_sdram_bankmachine4_cmd_payload_a <= videosoc_sdram_bankmachine4_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine4_cmd_payload_a <= {videosoc_sdram_bankmachine4_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine4_wait = (~((videosoc_sdram_bankmachine4_cmd_valid & videosoc_sdram_bankmachine4_cmd_ready) & videosoc_sdram_bankmachine4_cmd_payload_is_write));
assign videosoc_sdram_bankmachine4_syncfifo4_din = {videosoc_sdram_bankmachine4_fifo_in_last, videosoc_sdram_bankmachine4_fifo_in_first, videosoc_sdram_bankmachine4_fifo_in_payload_adr, videosoc_sdram_bankmachine4_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine4_fifo_out_last, videosoc_sdram_bankmachine4_fifo_out_first, videosoc_sdram_bankmachine4_fifo_out_payload_adr, videosoc_sdram_bankmachine4_fifo_out_payload_we} = videosoc_sdram_bankmachine4_syncfifo4_dout;
assign videosoc_sdram_bankmachine4_sink_ready = videosoc_sdram_bankmachine4_syncfifo4_writable;
assign videosoc_sdram_bankmachine4_syncfifo4_we = videosoc_sdram_bankmachine4_sink_valid;
assign videosoc_sdram_bankmachine4_fifo_in_first = videosoc_sdram_bankmachine4_sink_first;
assign videosoc_sdram_bankmachine4_fifo_in_last = videosoc_sdram_bankmachine4_sink_last;
assign videosoc_sdram_bankmachine4_fifo_in_payload_we = videosoc_sdram_bankmachine4_sink_payload_we;
assign videosoc_sdram_bankmachine4_fifo_in_payload_adr = videosoc_sdram_bankmachine4_sink_payload_adr;
assign videosoc_sdram_bankmachine4_source_valid = videosoc_sdram_bankmachine4_syncfifo4_readable;
assign videosoc_sdram_bankmachine4_source_first = videosoc_sdram_bankmachine4_fifo_out_first;
assign videosoc_sdram_bankmachine4_source_last = videosoc_sdram_bankmachine4_fifo_out_last;
assign videosoc_sdram_bankmachine4_source_payload_we = videosoc_sdram_bankmachine4_fifo_out_payload_we;
assign videosoc_sdram_bankmachine4_source_payload_adr = videosoc_sdram_bankmachine4_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine4_syncfifo4_re = videosoc_sdram_bankmachine4_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine4_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine4_replace) begin
		videosoc_sdram_bankmachine4_wrport_adr <= (videosoc_sdram_bankmachine4_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine4_wrport_adr <= videosoc_sdram_bankmachine4_produce;
	end
end
assign videosoc_sdram_bankmachine4_wrport_dat_w = videosoc_sdram_bankmachine4_syncfifo4_din;
assign videosoc_sdram_bankmachine4_wrport_we = (videosoc_sdram_bankmachine4_syncfifo4_we & (videosoc_sdram_bankmachine4_syncfifo4_writable | videosoc_sdram_bankmachine4_replace));
assign videosoc_sdram_bankmachine4_do_read = (videosoc_sdram_bankmachine4_syncfifo4_readable & videosoc_sdram_bankmachine4_syncfifo4_re);
assign videosoc_sdram_bankmachine4_rdport_adr = videosoc_sdram_bankmachine4_consume;
assign videosoc_sdram_bankmachine4_syncfifo4_dout = videosoc_sdram_bankmachine4_rdport_dat_r;
assign videosoc_sdram_bankmachine4_syncfifo4_writable = (videosoc_sdram_bankmachine4_level != 4'd8);
assign videosoc_sdram_bankmachine4_syncfifo4_readable = (videosoc_sdram_bankmachine4_level != 1'd0);
assign videosoc_sdram_bankmachine4_done = (videosoc_sdram_bankmachine4_count == 1'd0);
always @(*) begin
	videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd0;
	videosoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine4_req_wdata_ready <= 1'd0;
	bankmachine4_next_state <= 3'd0;
	videosoc_sdram_bankmachine4_req_rdata_valid <= 1'd0;
	videosoc_sdram_bankmachine4_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine4_cmd_valid <= 1'd0;
	videosoc_sdram_bankmachine4_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine4_track_open <= 1'd0;
	videosoc_sdram_bankmachine4_track_close <= 1'd0;
	videosoc_sdram_bankmachine4_cmd_payload_ras <= 1'd0;
	videosoc_sdram_bankmachine4_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine4_sel_row_adr <= 1'd0;
	bankmachine4_next_state <= bankmachine4_state;
	case (bankmachine4_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine4_done) begin
				videosoc_sdram_bankmachine4_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine4_cmd_ready) begin
					bankmachine4_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine4_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine4_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine4_track_open <= 1'd1;
			videosoc_sdram_bankmachine4_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine4_cmd_ready) begin
				bankmachine4_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine4_done) begin
				videosoc_sdram_bankmachine4_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine4_track_close <= 1'd1;
			videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine4_refresh_req)) begin
				bankmachine4_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine4_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine4_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine4_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine4_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine4_refresh_req) begin
				bankmachine4_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine4_source_valid) begin
					if (videosoc_sdram_bankmachine4_has_openrow) begin
						if (videosoc_sdram_bankmachine4_hit) begin
							videosoc_sdram_bankmachine4_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine4_source_payload_we) begin
								videosoc_sdram_bankmachine4_req_wdata_ready <= videosoc_sdram_bankmachine4_cmd_ready;
								videosoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine4_req_rdata_valid <= videosoc_sdram_bankmachine4_cmd_ready;
								videosoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine4_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine4_next_state <= 1'd1;
						end
					end else begin
						bankmachine4_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine5_sink_valid = videosoc_sdram_bankmachine5_req_valid;
assign videosoc_sdram_bankmachine5_req_ready = videosoc_sdram_bankmachine5_sink_ready;
assign videosoc_sdram_bankmachine5_sink_payload_we = videosoc_sdram_bankmachine5_req_we;
assign videosoc_sdram_bankmachine5_sink_payload_adr = videosoc_sdram_bankmachine5_req_adr;
assign videosoc_sdram_bankmachine5_source_ready = (videosoc_sdram_bankmachine5_req_wdata_ready | videosoc_sdram_bankmachine5_req_rdata_valid);
assign videosoc_sdram_bankmachine5_req_lock = videosoc_sdram_bankmachine5_source_valid;
assign videosoc_sdram_bankmachine5_hit = (videosoc_sdram_bankmachine5_openrow == videosoc_sdram_bankmachine5_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine5_cmd_payload_ba = 3'd5;
always @(*) begin
	videosoc_sdram_bankmachine5_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine5_sel_row_adr) begin
		videosoc_sdram_bankmachine5_cmd_payload_a <= videosoc_sdram_bankmachine5_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine5_cmd_payload_a <= {videosoc_sdram_bankmachine5_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine5_wait = (~((videosoc_sdram_bankmachine5_cmd_valid & videosoc_sdram_bankmachine5_cmd_ready) & videosoc_sdram_bankmachine5_cmd_payload_is_write));
assign videosoc_sdram_bankmachine5_syncfifo5_din = {videosoc_sdram_bankmachine5_fifo_in_last, videosoc_sdram_bankmachine5_fifo_in_first, videosoc_sdram_bankmachine5_fifo_in_payload_adr, videosoc_sdram_bankmachine5_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine5_fifo_out_last, videosoc_sdram_bankmachine5_fifo_out_first, videosoc_sdram_bankmachine5_fifo_out_payload_adr, videosoc_sdram_bankmachine5_fifo_out_payload_we} = videosoc_sdram_bankmachine5_syncfifo5_dout;
assign videosoc_sdram_bankmachine5_sink_ready = videosoc_sdram_bankmachine5_syncfifo5_writable;
assign videosoc_sdram_bankmachine5_syncfifo5_we = videosoc_sdram_bankmachine5_sink_valid;
assign videosoc_sdram_bankmachine5_fifo_in_first = videosoc_sdram_bankmachine5_sink_first;
assign videosoc_sdram_bankmachine5_fifo_in_last = videosoc_sdram_bankmachine5_sink_last;
assign videosoc_sdram_bankmachine5_fifo_in_payload_we = videosoc_sdram_bankmachine5_sink_payload_we;
assign videosoc_sdram_bankmachine5_fifo_in_payload_adr = videosoc_sdram_bankmachine5_sink_payload_adr;
assign videosoc_sdram_bankmachine5_source_valid = videosoc_sdram_bankmachine5_syncfifo5_readable;
assign videosoc_sdram_bankmachine5_source_first = videosoc_sdram_bankmachine5_fifo_out_first;
assign videosoc_sdram_bankmachine5_source_last = videosoc_sdram_bankmachine5_fifo_out_last;
assign videosoc_sdram_bankmachine5_source_payload_we = videosoc_sdram_bankmachine5_fifo_out_payload_we;
assign videosoc_sdram_bankmachine5_source_payload_adr = videosoc_sdram_bankmachine5_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine5_syncfifo5_re = videosoc_sdram_bankmachine5_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine5_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine5_replace) begin
		videosoc_sdram_bankmachine5_wrport_adr <= (videosoc_sdram_bankmachine5_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine5_wrport_adr <= videosoc_sdram_bankmachine5_produce;
	end
end
assign videosoc_sdram_bankmachine5_wrport_dat_w = videosoc_sdram_bankmachine5_syncfifo5_din;
assign videosoc_sdram_bankmachine5_wrport_we = (videosoc_sdram_bankmachine5_syncfifo5_we & (videosoc_sdram_bankmachine5_syncfifo5_writable | videosoc_sdram_bankmachine5_replace));
assign videosoc_sdram_bankmachine5_do_read = (videosoc_sdram_bankmachine5_syncfifo5_readable & videosoc_sdram_bankmachine5_syncfifo5_re);
assign videosoc_sdram_bankmachine5_rdport_adr = videosoc_sdram_bankmachine5_consume;
assign videosoc_sdram_bankmachine5_syncfifo5_dout = videosoc_sdram_bankmachine5_rdport_dat_r;
assign videosoc_sdram_bankmachine5_syncfifo5_writable = (videosoc_sdram_bankmachine5_level != 4'd8);
assign videosoc_sdram_bankmachine5_syncfifo5_readable = (videosoc_sdram_bankmachine5_level != 1'd0);
assign videosoc_sdram_bankmachine5_done = (videosoc_sdram_bankmachine5_count == 1'd0);
always @(*) begin
	bankmachine5_next_state <= 3'd0;
	videosoc_sdram_bankmachine5_track_open <= 1'd0;
	videosoc_sdram_bankmachine5_track_close <= 1'd0;
	videosoc_sdram_bankmachine5_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine5_cmd_payload_ras <= 1'd0;
	videosoc_sdram_bankmachine5_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine5_sel_row_adr <= 1'd0;
	videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd0;
	videosoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine5_req_wdata_ready <= 1'd0;
	videosoc_sdram_bankmachine5_req_rdata_valid <= 1'd0;
	videosoc_sdram_bankmachine5_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine5_cmd_valid <= 1'd0;
	bankmachine5_next_state <= bankmachine5_state;
	case (bankmachine5_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine5_done) begin
				videosoc_sdram_bankmachine5_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine5_cmd_ready) begin
					bankmachine5_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine5_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine5_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine5_track_open <= 1'd1;
			videosoc_sdram_bankmachine5_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine5_cmd_ready) begin
				bankmachine5_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine5_done) begin
				videosoc_sdram_bankmachine5_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine5_track_close <= 1'd1;
			videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine5_refresh_req)) begin
				bankmachine5_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine5_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine5_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine5_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine5_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine5_refresh_req) begin
				bankmachine5_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine5_source_valid) begin
					if (videosoc_sdram_bankmachine5_has_openrow) begin
						if (videosoc_sdram_bankmachine5_hit) begin
							videosoc_sdram_bankmachine5_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine5_source_payload_we) begin
								videosoc_sdram_bankmachine5_req_wdata_ready <= videosoc_sdram_bankmachine5_cmd_ready;
								videosoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine5_req_rdata_valid <= videosoc_sdram_bankmachine5_cmd_ready;
								videosoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine5_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine5_next_state <= 1'd1;
						end
					end else begin
						bankmachine5_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine6_sink_valid = videosoc_sdram_bankmachine6_req_valid;
assign videosoc_sdram_bankmachine6_req_ready = videosoc_sdram_bankmachine6_sink_ready;
assign videosoc_sdram_bankmachine6_sink_payload_we = videosoc_sdram_bankmachine6_req_we;
assign videosoc_sdram_bankmachine6_sink_payload_adr = videosoc_sdram_bankmachine6_req_adr;
assign videosoc_sdram_bankmachine6_source_ready = (videosoc_sdram_bankmachine6_req_wdata_ready | videosoc_sdram_bankmachine6_req_rdata_valid);
assign videosoc_sdram_bankmachine6_req_lock = videosoc_sdram_bankmachine6_source_valid;
assign videosoc_sdram_bankmachine6_hit = (videosoc_sdram_bankmachine6_openrow == videosoc_sdram_bankmachine6_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine6_cmd_payload_ba = 3'd6;
always @(*) begin
	videosoc_sdram_bankmachine6_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine6_sel_row_adr) begin
		videosoc_sdram_bankmachine6_cmd_payload_a <= videosoc_sdram_bankmachine6_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine6_cmd_payload_a <= {videosoc_sdram_bankmachine6_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine6_wait = (~((videosoc_sdram_bankmachine6_cmd_valid & videosoc_sdram_bankmachine6_cmd_ready) & videosoc_sdram_bankmachine6_cmd_payload_is_write));
assign videosoc_sdram_bankmachine6_syncfifo6_din = {videosoc_sdram_bankmachine6_fifo_in_last, videosoc_sdram_bankmachine6_fifo_in_first, videosoc_sdram_bankmachine6_fifo_in_payload_adr, videosoc_sdram_bankmachine6_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine6_fifo_out_last, videosoc_sdram_bankmachine6_fifo_out_first, videosoc_sdram_bankmachine6_fifo_out_payload_adr, videosoc_sdram_bankmachine6_fifo_out_payload_we} = videosoc_sdram_bankmachine6_syncfifo6_dout;
assign videosoc_sdram_bankmachine6_sink_ready = videosoc_sdram_bankmachine6_syncfifo6_writable;
assign videosoc_sdram_bankmachine6_syncfifo6_we = videosoc_sdram_bankmachine6_sink_valid;
assign videosoc_sdram_bankmachine6_fifo_in_first = videosoc_sdram_bankmachine6_sink_first;
assign videosoc_sdram_bankmachine6_fifo_in_last = videosoc_sdram_bankmachine6_sink_last;
assign videosoc_sdram_bankmachine6_fifo_in_payload_we = videosoc_sdram_bankmachine6_sink_payload_we;
assign videosoc_sdram_bankmachine6_fifo_in_payload_adr = videosoc_sdram_bankmachine6_sink_payload_adr;
assign videosoc_sdram_bankmachine6_source_valid = videosoc_sdram_bankmachine6_syncfifo6_readable;
assign videosoc_sdram_bankmachine6_source_first = videosoc_sdram_bankmachine6_fifo_out_first;
assign videosoc_sdram_bankmachine6_source_last = videosoc_sdram_bankmachine6_fifo_out_last;
assign videosoc_sdram_bankmachine6_source_payload_we = videosoc_sdram_bankmachine6_fifo_out_payload_we;
assign videosoc_sdram_bankmachine6_source_payload_adr = videosoc_sdram_bankmachine6_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine6_syncfifo6_re = videosoc_sdram_bankmachine6_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine6_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine6_replace) begin
		videosoc_sdram_bankmachine6_wrport_adr <= (videosoc_sdram_bankmachine6_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine6_wrport_adr <= videosoc_sdram_bankmachine6_produce;
	end
end
assign videosoc_sdram_bankmachine6_wrport_dat_w = videosoc_sdram_bankmachine6_syncfifo6_din;
assign videosoc_sdram_bankmachine6_wrport_we = (videosoc_sdram_bankmachine6_syncfifo6_we & (videosoc_sdram_bankmachine6_syncfifo6_writable | videosoc_sdram_bankmachine6_replace));
assign videosoc_sdram_bankmachine6_do_read = (videosoc_sdram_bankmachine6_syncfifo6_readable & videosoc_sdram_bankmachine6_syncfifo6_re);
assign videosoc_sdram_bankmachine6_rdport_adr = videosoc_sdram_bankmachine6_consume;
assign videosoc_sdram_bankmachine6_syncfifo6_dout = videosoc_sdram_bankmachine6_rdport_dat_r;
assign videosoc_sdram_bankmachine6_syncfifo6_writable = (videosoc_sdram_bankmachine6_level != 4'd8);
assign videosoc_sdram_bankmachine6_syncfifo6_readable = (videosoc_sdram_bankmachine6_level != 1'd0);
assign videosoc_sdram_bankmachine6_done = (videosoc_sdram_bankmachine6_count == 1'd0);
always @(*) begin
	videosoc_sdram_bankmachine6_req_rdata_valid <= 1'd0;
	videosoc_sdram_bankmachine6_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine6_cmd_valid <= 1'd0;
	videosoc_sdram_bankmachine6_track_open <= 1'd0;
	videosoc_sdram_bankmachine6_track_close <= 1'd0;
	videosoc_sdram_bankmachine6_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine6_cmd_payload_ras <= 1'd0;
	videosoc_sdram_bankmachine6_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine6_sel_row_adr <= 1'd0;
	videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd0;
	bankmachine6_next_state <= 3'd0;
	videosoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine6_req_wdata_ready <= 1'd0;
	bankmachine6_next_state <= bankmachine6_state;
	case (bankmachine6_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine6_done) begin
				videosoc_sdram_bankmachine6_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine6_cmd_ready) begin
					bankmachine6_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine6_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine6_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine6_track_open <= 1'd1;
			videosoc_sdram_bankmachine6_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine6_cmd_ready) begin
				bankmachine6_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine6_done) begin
				videosoc_sdram_bankmachine6_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine6_track_close <= 1'd1;
			videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine6_refresh_req)) begin
				bankmachine6_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine6_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine6_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine6_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine6_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine6_refresh_req) begin
				bankmachine6_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine6_source_valid) begin
					if (videosoc_sdram_bankmachine6_has_openrow) begin
						if (videosoc_sdram_bankmachine6_hit) begin
							videosoc_sdram_bankmachine6_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine6_source_payload_we) begin
								videosoc_sdram_bankmachine6_req_wdata_ready <= videosoc_sdram_bankmachine6_cmd_ready;
								videosoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine6_req_rdata_valid <= videosoc_sdram_bankmachine6_cmd_ready;
								videosoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine6_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine6_next_state <= 1'd1;
						end
					end else begin
						bankmachine6_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_bankmachine7_sink_valid = videosoc_sdram_bankmachine7_req_valid;
assign videosoc_sdram_bankmachine7_req_ready = videosoc_sdram_bankmachine7_sink_ready;
assign videosoc_sdram_bankmachine7_sink_payload_we = videosoc_sdram_bankmachine7_req_we;
assign videosoc_sdram_bankmachine7_sink_payload_adr = videosoc_sdram_bankmachine7_req_adr;
assign videosoc_sdram_bankmachine7_source_ready = (videosoc_sdram_bankmachine7_req_wdata_ready | videosoc_sdram_bankmachine7_req_rdata_valid);
assign videosoc_sdram_bankmachine7_req_lock = videosoc_sdram_bankmachine7_source_valid;
assign videosoc_sdram_bankmachine7_hit = (videosoc_sdram_bankmachine7_openrow == videosoc_sdram_bankmachine7_source_payload_adr[21:7]);
assign videosoc_sdram_bankmachine7_cmd_payload_ba = 3'd7;
always @(*) begin
	videosoc_sdram_bankmachine7_cmd_payload_a <= 15'd0;
	if (videosoc_sdram_bankmachine7_sel_row_adr) begin
		videosoc_sdram_bankmachine7_cmd_payload_a <= videosoc_sdram_bankmachine7_source_payload_adr[21:7];
	end else begin
		videosoc_sdram_bankmachine7_cmd_payload_a <= {videosoc_sdram_bankmachine7_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign videosoc_sdram_bankmachine7_wait = (~((videosoc_sdram_bankmachine7_cmd_valid & videosoc_sdram_bankmachine7_cmd_ready) & videosoc_sdram_bankmachine7_cmd_payload_is_write));
assign videosoc_sdram_bankmachine7_syncfifo7_din = {videosoc_sdram_bankmachine7_fifo_in_last, videosoc_sdram_bankmachine7_fifo_in_first, videosoc_sdram_bankmachine7_fifo_in_payload_adr, videosoc_sdram_bankmachine7_fifo_in_payload_we};
assign {videosoc_sdram_bankmachine7_fifo_out_last, videosoc_sdram_bankmachine7_fifo_out_first, videosoc_sdram_bankmachine7_fifo_out_payload_adr, videosoc_sdram_bankmachine7_fifo_out_payload_we} = videosoc_sdram_bankmachine7_syncfifo7_dout;
assign videosoc_sdram_bankmachine7_sink_ready = videosoc_sdram_bankmachine7_syncfifo7_writable;
assign videosoc_sdram_bankmachine7_syncfifo7_we = videosoc_sdram_bankmachine7_sink_valid;
assign videosoc_sdram_bankmachine7_fifo_in_first = videosoc_sdram_bankmachine7_sink_first;
assign videosoc_sdram_bankmachine7_fifo_in_last = videosoc_sdram_bankmachine7_sink_last;
assign videosoc_sdram_bankmachine7_fifo_in_payload_we = videosoc_sdram_bankmachine7_sink_payload_we;
assign videosoc_sdram_bankmachine7_fifo_in_payload_adr = videosoc_sdram_bankmachine7_sink_payload_adr;
assign videosoc_sdram_bankmachine7_source_valid = videosoc_sdram_bankmachine7_syncfifo7_readable;
assign videosoc_sdram_bankmachine7_source_first = videosoc_sdram_bankmachine7_fifo_out_first;
assign videosoc_sdram_bankmachine7_source_last = videosoc_sdram_bankmachine7_fifo_out_last;
assign videosoc_sdram_bankmachine7_source_payload_we = videosoc_sdram_bankmachine7_fifo_out_payload_we;
assign videosoc_sdram_bankmachine7_source_payload_adr = videosoc_sdram_bankmachine7_fifo_out_payload_adr;
assign videosoc_sdram_bankmachine7_syncfifo7_re = videosoc_sdram_bankmachine7_source_ready;
always @(*) begin
	videosoc_sdram_bankmachine7_wrport_adr <= 3'd0;
	if (videosoc_sdram_bankmachine7_replace) begin
		videosoc_sdram_bankmachine7_wrport_adr <= (videosoc_sdram_bankmachine7_produce - 1'd1);
	end else begin
		videosoc_sdram_bankmachine7_wrport_adr <= videosoc_sdram_bankmachine7_produce;
	end
end
assign videosoc_sdram_bankmachine7_wrport_dat_w = videosoc_sdram_bankmachine7_syncfifo7_din;
assign videosoc_sdram_bankmachine7_wrport_we = (videosoc_sdram_bankmachine7_syncfifo7_we & (videosoc_sdram_bankmachine7_syncfifo7_writable | videosoc_sdram_bankmachine7_replace));
assign videosoc_sdram_bankmachine7_do_read = (videosoc_sdram_bankmachine7_syncfifo7_readable & videosoc_sdram_bankmachine7_syncfifo7_re);
assign videosoc_sdram_bankmachine7_rdport_adr = videosoc_sdram_bankmachine7_consume;
assign videosoc_sdram_bankmachine7_syncfifo7_dout = videosoc_sdram_bankmachine7_rdport_dat_r;
assign videosoc_sdram_bankmachine7_syncfifo7_writable = (videosoc_sdram_bankmachine7_level != 4'd8);
assign videosoc_sdram_bankmachine7_syncfifo7_readable = (videosoc_sdram_bankmachine7_level != 1'd0);
assign videosoc_sdram_bankmachine7_done = (videosoc_sdram_bankmachine7_count == 1'd0);
always @(*) begin
	videosoc_sdram_bankmachine7_cmd_payload_ras <= 1'd0;
	videosoc_sdram_bankmachine7_cmd_payload_we <= 1'd0;
	videosoc_sdram_bankmachine7_sel_row_adr <= 1'd0;
	videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd0;
	videosoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd0;
	videosoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd0;
	videosoc_sdram_bankmachine7_req_wdata_ready <= 1'd0;
	videosoc_sdram_bankmachine7_req_rdata_valid <= 1'd0;
	videosoc_sdram_bankmachine7_refresh_gnt <= 1'd0;
	videosoc_sdram_bankmachine7_cmd_valid <= 1'd0;
	bankmachine7_next_state <= 3'd0;
	videosoc_sdram_bankmachine7_cmd_payload_cas <= 1'd0;
	videosoc_sdram_bankmachine7_track_open <= 1'd0;
	videosoc_sdram_bankmachine7_track_close <= 1'd0;
	bankmachine7_next_state <= bankmachine7_state;
	case (bankmachine7_state)
		1'd1: begin
			if (videosoc_sdram_bankmachine7_done) begin
				videosoc_sdram_bankmachine7_cmd_valid <= 1'd1;
				if (videosoc_sdram_bankmachine7_cmd_ready) begin
					bankmachine7_next_state <= 3'd4;
				end
				videosoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
				videosoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
				videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			end
			videosoc_sdram_bankmachine7_track_close <= 1'd1;
		end
		2'd2: begin
			videosoc_sdram_bankmachine7_sel_row_adr <= 1'd1;
			videosoc_sdram_bankmachine7_track_open <= 1'd1;
			videosoc_sdram_bankmachine7_cmd_valid <= 1'd1;
			videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if (videosoc_sdram_bankmachine7_cmd_ready) begin
				bankmachine7_next_state <= 3'd6;
			end
			videosoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (videosoc_sdram_bankmachine7_done) begin
				videosoc_sdram_bankmachine7_refresh_gnt <= 1'd1;
			end
			videosoc_sdram_bankmachine7_track_close <= 1'd1;
			videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if ((~videosoc_sdram_bankmachine7_refresh_req)) begin
				bankmachine7_next_state <= 1'd0;
			end
		end
		3'd4: begin
			bankmachine7_next_state <= 3'd5;
		end
		3'd5: begin
			bankmachine7_next_state <= 2'd2;
		end
		3'd6: begin
			bankmachine7_next_state <= 3'd7;
		end
		3'd7: begin
			bankmachine7_next_state <= 1'd0;
		end
		default: begin
			if (videosoc_sdram_bankmachine7_refresh_req) begin
				bankmachine7_next_state <= 2'd3;
			end else begin
				if (videosoc_sdram_bankmachine7_source_valid) begin
					if (videosoc_sdram_bankmachine7_has_openrow) begin
						if (videosoc_sdram_bankmachine7_hit) begin
							videosoc_sdram_bankmachine7_cmd_valid <= 1'd1;
							if (videosoc_sdram_bankmachine7_source_payload_we) begin
								videosoc_sdram_bankmachine7_req_wdata_ready <= videosoc_sdram_bankmachine7_cmd_ready;
								videosoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd1;
								videosoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
							end else begin
								videosoc_sdram_bankmachine7_req_rdata_valid <= videosoc_sdram_bankmachine7_cmd_ready;
								videosoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd1;
							end
							videosoc_sdram_bankmachine7_cmd_payload_cas <= 1'd1;
						end else begin
							bankmachine7_next_state <= 1'd1;
						end
					end else begin
						bankmachine7_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign videosoc_sdram_read_available = ((((((((videosoc_sdram_bankmachine0_cmd_valid & videosoc_sdram_bankmachine0_cmd_payload_is_read) | (videosoc_sdram_bankmachine1_cmd_valid & videosoc_sdram_bankmachine1_cmd_payload_is_read)) | (videosoc_sdram_bankmachine2_cmd_valid & videosoc_sdram_bankmachine2_cmd_payload_is_read)) | (videosoc_sdram_bankmachine3_cmd_valid & videosoc_sdram_bankmachine3_cmd_payload_is_read)) | (videosoc_sdram_bankmachine4_cmd_valid & videosoc_sdram_bankmachine4_cmd_payload_is_read)) | (videosoc_sdram_bankmachine5_cmd_valid & videosoc_sdram_bankmachine5_cmd_payload_is_read)) | (videosoc_sdram_bankmachine6_cmd_valid & videosoc_sdram_bankmachine6_cmd_payload_is_read)) | (videosoc_sdram_bankmachine7_cmd_valid & videosoc_sdram_bankmachine7_cmd_payload_is_read));
assign videosoc_sdram_write_available = ((((((((videosoc_sdram_bankmachine0_cmd_valid & videosoc_sdram_bankmachine0_cmd_payload_is_write) | (videosoc_sdram_bankmachine1_cmd_valid & videosoc_sdram_bankmachine1_cmd_payload_is_write)) | (videosoc_sdram_bankmachine2_cmd_valid & videosoc_sdram_bankmachine2_cmd_payload_is_write)) | (videosoc_sdram_bankmachine3_cmd_valid & videosoc_sdram_bankmachine3_cmd_payload_is_write)) | (videosoc_sdram_bankmachine4_cmd_valid & videosoc_sdram_bankmachine4_cmd_payload_is_write)) | (videosoc_sdram_bankmachine5_cmd_valid & videosoc_sdram_bankmachine5_cmd_payload_is_write)) | (videosoc_sdram_bankmachine6_cmd_valid & videosoc_sdram_bankmachine6_cmd_payload_is_write)) | (videosoc_sdram_bankmachine7_cmd_valid & videosoc_sdram_bankmachine7_cmd_payload_is_write));
assign videosoc_sdram_max_time0 = (videosoc_sdram_time0 == 1'd0);
assign videosoc_sdram_max_time1 = (videosoc_sdram_time1 == 1'd0);
assign videosoc_sdram_bankmachine0_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_bankmachine1_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_bankmachine2_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_bankmachine3_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_bankmachine4_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_bankmachine5_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_bankmachine6_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_bankmachine7_refresh_req = videosoc_sdram_cmd_valid;
assign videosoc_sdram_go_to_refresh = (((((((videosoc_sdram_bankmachine0_refresh_gnt & videosoc_sdram_bankmachine1_refresh_gnt) & videosoc_sdram_bankmachine2_refresh_gnt) & videosoc_sdram_bankmachine3_refresh_gnt) & videosoc_sdram_bankmachine4_refresh_gnt) & videosoc_sdram_bankmachine5_refresh_gnt) & videosoc_sdram_bankmachine6_refresh_gnt) & videosoc_sdram_bankmachine7_refresh_gnt);
assign videosoc_sdram_interface_rdata = {videosoc_sdram_dfi_p3_rddata, videosoc_sdram_dfi_p2_rddata, videosoc_sdram_dfi_p1_rddata, videosoc_sdram_dfi_p0_rddata};
assign {videosoc_sdram_dfi_p3_wrdata, videosoc_sdram_dfi_p2_wrdata, videosoc_sdram_dfi_p1_wrdata, videosoc_sdram_dfi_p0_wrdata} = videosoc_sdram_interface_wdata;
assign {videosoc_sdram_dfi_p3_wrdata_mask, videosoc_sdram_dfi_p2_wrdata_mask, videosoc_sdram_dfi_p1_wrdata_mask, videosoc_sdram_dfi_p0_wrdata_mask} = (~videosoc_sdram_interface_wdata_we);
always @(*) begin
	videosoc_sdram_choose_cmd_valids <= 8'd0;
	videosoc_sdram_choose_cmd_valids[0] <= (videosoc_sdram_bankmachine0_cmd_valid & ((videosoc_sdram_bankmachine0_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine0_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine0_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
	videosoc_sdram_choose_cmd_valids[1] <= (videosoc_sdram_bankmachine1_cmd_valid & ((videosoc_sdram_bankmachine1_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine1_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine1_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
	videosoc_sdram_choose_cmd_valids[2] <= (videosoc_sdram_bankmachine2_cmd_valid & ((videosoc_sdram_bankmachine2_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine2_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine2_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
	videosoc_sdram_choose_cmd_valids[3] <= (videosoc_sdram_bankmachine3_cmd_valid & ((videosoc_sdram_bankmachine3_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine3_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine3_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
	videosoc_sdram_choose_cmd_valids[4] <= (videosoc_sdram_bankmachine4_cmd_valid & ((videosoc_sdram_bankmachine4_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine4_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine4_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
	videosoc_sdram_choose_cmd_valids[5] <= (videosoc_sdram_bankmachine5_cmd_valid & ((videosoc_sdram_bankmachine5_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine5_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine5_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
	videosoc_sdram_choose_cmd_valids[6] <= (videosoc_sdram_bankmachine6_cmd_valid & ((videosoc_sdram_bankmachine6_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine6_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine6_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
	videosoc_sdram_choose_cmd_valids[7] <= (videosoc_sdram_bankmachine7_cmd_valid & ((videosoc_sdram_bankmachine7_cmd_payload_is_cmd & videosoc_sdram_choose_cmd_want_cmds) | ((videosoc_sdram_bankmachine7_cmd_payload_is_read == videosoc_sdram_choose_cmd_want_reads) & (videosoc_sdram_bankmachine7_cmd_payload_is_write == videosoc_sdram_choose_cmd_want_writes))));
end
assign videosoc_sdram_choose_cmd_request = videosoc_sdram_choose_cmd_valids;
assign videosoc_sdram_choose_cmd_cmd_valid = comb_rhs_array_muxed0;
assign videosoc_sdram_choose_cmd_cmd_payload_a = comb_rhs_array_muxed1;
assign videosoc_sdram_choose_cmd_cmd_payload_ba = comb_rhs_array_muxed2;
assign videosoc_sdram_choose_cmd_cmd_payload_is_read = comb_rhs_array_muxed3;
assign videosoc_sdram_choose_cmd_cmd_payload_is_write = comb_rhs_array_muxed4;
assign videosoc_sdram_choose_cmd_cmd_payload_is_cmd = comb_rhs_array_muxed5;
always @(*) begin
	videosoc_sdram_choose_cmd_cmd_payload_cas <= 1'd0;
	if (videosoc_sdram_choose_cmd_cmd_valid) begin
		videosoc_sdram_choose_cmd_cmd_payload_cas <= comb_t_array_muxed0;
	end
end
always @(*) begin
	videosoc_sdram_choose_cmd_cmd_payload_ras <= 1'd0;
	if (videosoc_sdram_choose_cmd_cmd_valid) begin
		videosoc_sdram_choose_cmd_cmd_payload_ras <= comb_t_array_muxed1;
	end
end
always @(*) begin
	videosoc_sdram_choose_cmd_cmd_payload_we <= 1'd0;
	if (videosoc_sdram_choose_cmd_cmd_valid) begin
		videosoc_sdram_choose_cmd_cmd_payload_we <= comb_t_array_muxed2;
	end
end
assign videosoc_sdram_choose_cmd_ce = videosoc_sdram_choose_cmd_cmd_ready;
always @(*) begin
	videosoc_sdram_choose_req_valids <= 8'd0;
	videosoc_sdram_choose_req_valids[0] <= (videosoc_sdram_bankmachine0_cmd_valid & ((videosoc_sdram_bankmachine0_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine0_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine0_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
	videosoc_sdram_choose_req_valids[1] <= (videosoc_sdram_bankmachine1_cmd_valid & ((videosoc_sdram_bankmachine1_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine1_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine1_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
	videosoc_sdram_choose_req_valids[2] <= (videosoc_sdram_bankmachine2_cmd_valid & ((videosoc_sdram_bankmachine2_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine2_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine2_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
	videosoc_sdram_choose_req_valids[3] <= (videosoc_sdram_bankmachine3_cmd_valid & ((videosoc_sdram_bankmachine3_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine3_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine3_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
	videosoc_sdram_choose_req_valids[4] <= (videosoc_sdram_bankmachine4_cmd_valid & ((videosoc_sdram_bankmachine4_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine4_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine4_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
	videosoc_sdram_choose_req_valids[5] <= (videosoc_sdram_bankmachine5_cmd_valid & ((videosoc_sdram_bankmachine5_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine5_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine5_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
	videosoc_sdram_choose_req_valids[6] <= (videosoc_sdram_bankmachine6_cmd_valid & ((videosoc_sdram_bankmachine6_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine6_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine6_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
	videosoc_sdram_choose_req_valids[7] <= (videosoc_sdram_bankmachine7_cmd_valid & ((videosoc_sdram_bankmachine7_cmd_payload_is_cmd & videosoc_sdram_choose_req_want_cmds) | ((videosoc_sdram_bankmachine7_cmd_payload_is_read == videosoc_sdram_choose_req_want_reads) & (videosoc_sdram_bankmachine7_cmd_payload_is_write == videosoc_sdram_choose_req_want_writes))));
end
assign videosoc_sdram_choose_req_request = videosoc_sdram_choose_req_valids;
assign videosoc_sdram_choose_req_cmd_valid = comb_rhs_array_muxed6;
assign videosoc_sdram_choose_req_cmd_payload_a = comb_rhs_array_muxed7;
assign videosoc_sdram_choose_req_cmd_payload_ba = comb_rhs_array_muxed8;
assign videosoc_sdram_choose_req_cmd_payload_is_read = comb_rhs_array_muxed9;
assign videosoc_sdram_choose_req_cmd_payload_is_write = comb_rhs_array_muxed10;
assign videosoc_sdram_choose_req_cmd_payload_is_cmd = comb_rhs_array_muxed11;
always @(*) begin
	videosoc_sdram_choose_req_cmd_payload_cas <= 1'd0;
	if (videosoc_sdram_choose_req_cmd_valid) begin
		videosoc_sdram_choose_req_cmd_payload_cas <= comb_t_array_muxed3;
	end
end
always @(*) begin
	videosoc_sdram_choose_req_cmd_payload_ras <= 1'd0;
	if (videosoc_sdram_choose_req_cmd_valid) begin
		videosoc_sdram_choose_req_cmd_payload_ras <= comb_t_array_muxed4;
	end
end
always @(*) begin
	videosoc_sdram_choose_req_cmd_payload_we <= 1'd0;
	if (videosoc_sdram_choose_req_cmd_valid) begin
		videosoc_sdram_choose_req_cmd_payload_we <= comb_t_array_muxed5;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine0_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 1'd0))) begin
		videosoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 1'd0))) begin
		videosoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine1_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 1'd1))) begin
		videosoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 1'd1))) begin
		videosoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine2_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 2'd2))) begin
		videosoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 2'd2))) begin
		videosoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine3_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 2'd3))) begin
		videosoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 2'd3))) begin
		videosoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine4_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 3'd4))) begin
		videosoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 3'd4))) begin
		videosoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine5_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 3'd5))) begin
		videosoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 3'd5))) begin
		videosoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine6_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 3'd6))) begin
		videosoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 3'd6))) begin
		videosoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	videosoc_sdram_bankmachine7_cmd_ready <= 1'd0;
	if (((videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_ready) & (videosoc_sdram_choose_cmd_grant == 3'd7))) begin
		videosoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
	if (((videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_ready) & (videosoc_sdram_choose_req_grant == 3'd7))) begin
		videosoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
end
assign videosoc_sdram_choose_req_ce = videosoc_sdram_choose_req_cmd_ready;
assign videosoc_sdram_dfi_p0_cke = 1'd1;
assign videosoc_sdram_dfi_p0_cs_n = 1'd0;
assign videosoc_sdram_dfi_p0_odt = 1'd1;
assign videosoc_sdram_dfi_p0_reset_n = 1'd1;
assign videosoc_sdram_dfi_p1_cke = 1'd1;
assign videosoc_sdram_dfi_p1_cs_n = 1'd0;
assign videosoc_sdram_dfi_p1_odt = 1'd1;
assign videosoc_sdram_dfi_p1_reset_n = 1'd1;
assign videosoc_sdram_dfi_p2_cke = 1'd1;
assign videosoc_sdram_dfi_p2_cs_n = 1'd0;
assign videosoc_sdram_dfi_p2_odt = 1'd1;
assign videosoc_sdram_dfi_p2_reset_n = 1'd1;
assign videosoc_sdram_dfi_p3_cke = 1'd1;
assign videosoc_sdram_dfi_p3_cs_n = 1'd0;
assign videosoc_sdram_dfi_p3_odt = 1'd1;
assign videosoc_sdram_dfi_p3_reset_n = 1'd1;
always @(*) begin
	videosoc_sdram_choose_req_cmd_ready <= 1'd0;
	videosoc_sdram_en1 <= 1'd0;
	videosoc_sdram_cmd_ready <= 1'd0;
	multiplexer_next_state <= 4'd0;
	videosoc_sdram_choose_cmd_cmd_ready <= 1'd0;
	videosoc_sdram_sel0 <= 2'd0;
	videosoc_sdram_sel1 <= 2'd0;
	videosoc_sdram_en0 <= 1'd0;
	videosoc_sdram_sel2 <= 2'd0;
	videosoc_sdram_sel3 <= 2'd0;
	videosoc_sdram_choose_req_want_reads <= 1'd0;
	videosoc_sdram_choose_req_want_writes <= 1'd0;
	multiplexer_next_state <= multiplexer_state;
	case (multiplexer_state)
		1'd1: begin
			videosoc_sdram_en1 <= 1'd1;
			videosoc_sdram_choose_req_want_writes <= 1'd1;
			videosoc_sdram_choose_cmd_cmd_ready <= 1'd1;
			videosoc_sdram_choose_req_cmd_ready <= 1'd1;
			videosoc_sdram_sel0 <= 1'd1;
			videosoc_sdram_sel1 <= 1'd0;
			videosoc_sdram_sel2 <= 2'd2;
			videosoc_sdram_sel3 <= 1'd0;
			if (videosoc_sdram_read_available) begin
				if (((~videosoc_sdram_write_available) | videosoc_sdram_max_time1)) begin
					multiplexer_next_state <= 4'd8;
				end
			end
			if (videosoc_sdram_go_to_refresh) begin
				multiplexer_next_state <= 2'd2;
			end
		end
		2'd2: begin
			videosoc_sdram_sel0 <= 2'd3;
			videosoc_sdram_cmd_ready <= 1'd1;
			if (videosoc_sdram_cmd_last) begin
				multiplexer_next_state <= 1'd0;
			end
		end
		2'd3: begin
			multiplexer_next_state <= 3'd4;
		end
		3'd4: begin
			multiplexer_next_state <= 3'd5;
		end
		3'd5: begin
			multiplexer_next_state <= 3'd6;
		end
		3'd6: begin
			multiplexer_next_state <= 3'd7;
		end
		3'd7: begin
			multiplexer_next_state <= 1'd1;
		end
		4'd8: begin
			multiplexer_next_state <= 4'd9;
		end
		4'd9: begin
			multiplexer_next_state <= 4'd10;
		end
		4'd10: begin
			multiplexer_next_state <= 4'd11;
		end
		4'd11: begin
			multiplexer_next_state <= 4'd12;
		end
		4'd12: begin
			multiplexer_next_state <= 4'd13;
		end
		4'd13: begin
			multiplexer_next_state <= 4'd14;
		end
		4'd14: begin
			multiplexer_next_state <= 1'd0;
		end
		default: begin
			videosoc_sdram_en0 <= 1'd1;
			videosoc_sdram_choose_req_want_reads <= 1'd1;
			videosoc_sdram_choose_cmd_cmd_ready <= 1'd1;
			videosoc_sdram_choose_req_cmd_ready <= 1'd1;
			videosoc_sdram_sel0 <= 2'd2;
			videosoc_sdram_sel1 <= 1'd1;
			videosoc_sdram_sel2 <= 1'd0;
			videosoc_sdram_sel3 <= 1'd0;
			if (videosoc_sdram_write_available) begin
				if (((~videosoc_sdram_read_available) | videosoc_sdram_max_time0)) begin
					multiplexer_next_state <= 2'd3;
				end
			end
			if (videosoc_sdram_go_to_refresh) begin
				multiplexer_next_state <= 2'd2;
			end
		end
	endcase
end
assign cba0 = videosoc_port_cmd_payload_adr[9:7];
assign rca0 = {videosoc_port_cmd_payload_adr[24:10], videosoc_port_cmd_payload_adr[6:0]};
assign cba1 = litedramcrossbar_cmd_payload_adr[9:7];
assign rca1 = {litedramcrossbar_cmd_payload_adr[24:10], litedramcrossbar_cmd_payload_adr[6:0]};
assign cba2 = hdmi_out0_dram_port_cmd_payload_adr[9:7];
assign rca2 = {hdmi_out0_dram_port_cmd_payload_adr[24:10], hdmi_out0_dram_port_cmd_payload_adr[6:0]};
assign roundrobin0_request = {(((cba2 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin0_ce = ((~videosoc_sdram_interface_bank0_valid) & (~videosoc_sdram_interface_bank0_lock));
assign videosoc_sdram_interface_bank0_adr = comb_rhs_array_muxed12;
assign videosoc_sdram_interface_bank0_we = comb_rhs_array_muxed13;
assign videosoc_sdram_interface_bank0_valid = comb_rhs_array_muxed14;
assign roundrobin1_request = {(((cba2 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin1_ce = ((~videosoc_sdram_interface_bank1_valid) & (~videosoc_sdram_interface_bank1_lock));
assign videosoc_sdram_interface_bank1_adr = comb_rhs_array_muxed15;
assign videosoc_sdram_interface_bank1_we = comb_rhs_array_muxed16;
assign videosoc_sdram_interface_bank1_valid = comb_rhs_array_muxed17;
assign roundrobin2_request = {(((cba2 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin2_ce = ((~videosoc_sdram_interface_bank2_valid) & (~videosoc_sdram_interface_bank2_lock));
assign videosoc_sdram_interface_bank2_adr = comb_rhs_array_muxed18;
assign videosoc_sdram_interface_bank2_we = comb_rhs_array_muxed19;
assign videosoc_sdram_interface_bank2_valid = comb_rhs_array_muxed20;
assign roundrobin3_request = {(((cba2 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin3_ce = ((~videosoc_sdram_interface_bank3_valid) & (~videosoc_sdram_interface_bank3_lock));
assign videosoc_sdram_interface_bank3_adr = comb_rhs_array_muxed21;
assign videosoc_sdram_interface_bank3_we = comb_rhs_array_muxed22;
assign videosoc_sdram_interface_bank3_valid = comb_rhs_array_muxed23;
assign roundrobin4_request = {(((cba2 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin4_ce = ((~videosoc_sdram_interface_bank4_valid) & (~videosoc_sdram_interface_bank4_lock));
assign videosoc_sdram_interface_bank4_adr = comb_rhs_array_muxed24;
assign videosoc_sdram_interface_bank4_we = comb_rhs_array_muxed25;
assign videosoc_sdram_interface_bank4_valid = comb_rhs_array_muxed26;
assign roundrobin5_request = {(((cba2 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin5_ce = ((~videosoc_sdram_interface_bank5_valid) & (~videosoc_sdram_interface_bank5_lock));
assign videosoc_sdram_interface_bank5_adr = comb_rhs_array_muxed27;
assign videosoc_sdram_interface_bank5_we = comb_rhs_array_muxed28;
assign videosoc_sdram_interface_bank5_valid = comb_rhs_array_muxed29;
assign roundrobin6_request = {(((cba2 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin6_ce = ((~videosoc_sdram_interface_bank6_valid) & (~videosoc_sdram_interface_bank6_lock));
assign videosoc_sdram_interface_bank6_adr = comb_rhs_array_muxed30;
assign videosoc_sdram_interface_bank6_we = comb_rhs_array_muxed31;
assign videosoc_sdram_interface_bank6_valid = comb_rhs_array_muxed32;
assign roundrobin7_request = {(((cba2 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid), (((cba1 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))))) & litedramcrossbar_cmd_valid), (((cba0 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))))) & videosoc_port_cmd_valid)};
assign roundrobin7_ce = ((~videosoc_sdram_interface_bank7_valid) & (~videosoc_sdram_interface_bank7_lock));
assign videosoc_sdram_interface_bank7_adr = comb_rhs_array_muxed33;
assign videosoc_sdram_interface_bank7_we = comb_rhs_array_muxed34;
assign videosoc_sdram_interface_bank7_valid = comb_rhs_array_muxed35;
assign videosoc_port_cmd_ready = ((((((((1'd0 | (((roundrobin0_grant == 1'd0) & ((cba0 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0)))))) & videosoc_sdram_interface_bank0_ready)) | (((roundrobin1_grant == 1'd0) & ((cba0 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0)))))) & videosoc_sdram_interface_bank1_ready)) | (((roundrobin2_grant == 1'd0) & ((cba0 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0)))))) & videosoc_sdram_interface_bank2_ready)) | (((roundrobin3_grant == 1'd0) & ((cba0 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0)))))) & videosoc_sdram_interface_bank3_ready)) | (((roundrobin4_grant == 1'd0) & ((cba0 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0)))))) & videosoc_sdram_interface_bank4_ready)) | (((roundrobin5_grant == 1'd0) & ((cba0 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0)))))) & videosoc_sdram_interface_bank5_ready)) | (((roundrobin6_grant == 1'd0) & ((cba0 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0)))))) & videosoc_sdram_interface_bank6_ready)) | (((roundrobin7_grant == 1'd0) & ((cba0 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0)))))) & videosoc_sdram_interface_bank7_ready));
assign litedramcrossbar_cmd_ready = ((((((((1'd0 | (((roundrobin0_grant == 1'd1) & ((cba1 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1)))))) & videosoc_sdram_interface_bank0_ready)) | (((roundrobin1_grant == 1'd1) & ((cba1 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1)))))) & videosoc_sdram_interface_bank1_ready)) | (((roundrobin2_grant == 1'd1) & ((cba1 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1)))))) & videosoc_sdram_interface_bank2_ready)) | (((roundrobin3_grant == 1'd1) & ((cba1 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1)))))) & videosoc_sdram_interface_bank3_ready)) | (((roundrobin4_grant == 1'd1) & ((cba1 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1)))))) & videosoc_sdram_interface_bank4_ready)) | (((roundrobin5_grant == 1'd1) & ((cba1 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1)))))) & videosoc_sdram_interface_bank5_ready)) | (((roundrobin6_grant == 1'd1) & ((cba1 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1)))))) & videosoc_sdram_interface_bank6_ready)) | (((roundrobin7_grant == 1'd1) & ((cba1 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1)))))) & videosoc_sdram_interface_bank7_ready));
assign hdmi_out0_dram_port_cmd_ready = ((((((((1'd0 | (((roundrobin0_grant == 2'd2) & ((cba2 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2)))))) & videosoc_sdram_interface_bank0_ready)) | (((roundrobin1_grant == 2'd2) & ((cba2 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2)))))) & videosoc_sdram_interface_bank1_ready)) | (((roundrobin2_grant == 2'd2) & ((cba2 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2)))))) & videosoc_sdram_interface_bank2_ready)) | (((roundrobin3_grant == 2'd2) & ((cba2 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2)))))) & videosoc_sdram_interface_bank3_ready)) | (((roundrobin4_grant == 2'd2) & ((cba2 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2)))))) & videosoc_sdram_interface_bank4_ready)) | (((roundrobin5_grant == 2'd2) & ((cba2 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2)))))) & videosoc_sdram_interface_bank5_ready)) | (((roundrobin6_grant == 2'd2) & ((cba2 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2)))))) & videosoc_sdram_interface_bank6_ready)) | (((roundrobin7_grant == 2'd2) & ((cba2 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2)))))) & videosoc_sdram_interface_bank7_ready));
assign videosoc_port_wdata_ready = new_master_wdata_ready2;
assign litedramcrossbar_wdata_ready = new_master_wdata_ready5;
assign hdmi_out0_dram_port_wdata_ready = new_master_wdata_ready8;
assign videosoc_port_rdata_valid = new_master_rdata_valid6;
assign litedramcrossbar_rdata_valid = new_master_rdata_valid13;
assign hdmi_out0_dram_port_rdata_valid = new_master_rdata_valid20;
always @(*) begin
	videosoc_sdram_interface_wdata <= 128'd0;
	videosoc_sdram_interface_wdata_we <= 16'd0;
	case ({new_master_wdata_ready8, new_master_wdata_ready5, new_master_wdata_ready2})
		1'd1: begin
			videosoc_sdram_interface_wdata <= videosoc_port_wdata_payload_data;
			videosoc_sdram_interface_wdata_we <= videosoc_port_wdata_payload_we;
		end
		2'd2: begin
			videosoc_sdram_interface_wdata <= litedramcrossbar_wdata_payload_data;
			videosoc_sdram_interface_wdata_we <= litedramcrossbar_wdata_payload_we;
		end
		3'd4: begin
			videosoc_sdram_interface_wdata <= hdmi_out0_dram_port_wdata_payload_data;
			videosoc_sdram_interface_wdata_we <= hdmi_out0_dram_port_wdata_payload_we;
		end
		default: begin
			videosoc_sdram_interface_wdata <= 1'd0;
			videosoc_sdram_interface_wdata_we <= 1'd0;
		end
	endcase
end
assign videosoc_port_rdata_payload_data = videosoc_sdram_interface_rdata;
assign litedramcrossbar_rdata_payload_data = videosoc_sdram_interface_rdata;
assign hdmi_out0_dram_port_rdata_payload_data = videosoc_sdram_interface_rdata;
assign hdmi_out0_dram_port_cmd_fifo_asyncfifo_din = {hdmi_out0_dram_port_cmd_fifo_fifo_in_last, hdmi_out0_dram_port_cmd_fifo_fifo_in_first, hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_adr, hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_we};
assign {hdmi_out0_dram_port_cmd_fifo_fifo_out_last, hdmi_out0_dram_port_cmd_fifo_fifo_out_first, hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_adr, hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_we} = hdmi_out0_dram_port_cmd_fifo_asyncfifo_dout;
assign hdmi_out0_dram_port_cmd_fifo_sink_ready = hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable;
assign hdmi_out0_dram_port_cmd_fifo_asyncfifo_we = hdmi_out0_dram_port_cmd_fifo_sink_valid;
assign hdmi_out0_dram_port_cmd_fifo_fifo_in_first = hdmi_out0_dram_port_cmd_fifo_sink_first;
assign hdmi_out0_dram_port_cmd_fifo_fifo_in_last = hdmi_out0_dram_port_cmd_fifo_sink_last;
assign hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_we = hdmi_out0_dram_port_cmd_fifo_sink_payload_we;
assign hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_adr = hdmi_out0_dram_port_cmd_fifo_sink_payload_adr;
assign hdmi_out0_dram_port_cmd_fifo_source_valid = hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable;
assign hdmi_out0_dram_port_cmd_fifo_source_first = hdmi_out0_dram_port_cmd_fifo_fifo_out_first;
assign hdmi_out0_dram_port_cmd_fifo_source_last = hdmi_out0_dram_port_cmd_fifo_fifo_out_last;
assign hdmi_out0_dram_port_cmd_fifo_source_payload_we = hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_we;
assign hdmi_out0_dram_port_cmd_fifo_source_payload_adr = hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_adr;
assign hdmi_out0_dram_port_cmd_fifo_asyncfifo_re = hdmi_out0_dram_port_cmd_fifo_source_ready;
assign hdmi_out0_dram_port_cmd_fifo_graycounter0_ce = (hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable & hdmi_out0_dram_port_cmd_fifo_asyncfifo_we);
assign hdmi_out0_dram_port_cmd_fifo_graycounter1_ce = (hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable & hdmi_out0_dram_port_cmd_fifo_asyncfifo_re);
assign hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable = (((hdmi_out0_dram_port_cmd_fifo_graycounter0_q[2] == hdmi_out0_dram_port_cmd_fifo_consume_wdomain[2]) | (hdmi_out0_dram_port_cmd_fifo_graycounter0_q[1] == hdmi_out0_dram_port_cmd_fifo_consume_wdomain[1])) | (hdmi_out0_dram_port_cmd_fifo_graycounter0_q[0] != hdmi_out0_dram_port_cmd_fifo_consume_wdomain[0]));
assign hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable = (hdmi_out0_dram_port_cmd_fifo_graycounter1_q != hdmi_out0_dram_port_cmd_fifo_produce_rdomain);
assign hdmi_out0_dram_port_cmd_fifo_wrport_adr = hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary[1:0];
assign hdmi_out0_dram_port_cmd_fifo_wrport_dat_w = hdmi_out0_dram_port_cmd_fifo_asyncfifo_din;
assign hdmi_out0_dram_port_cmd_fifo_wrport_we = hdmi_out0_dram_port_cmd_fifo_graycounter0_ce;
assign hdmi_out0_dram_port_cmd_fifo_rdport_adr = hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary[1:0];
assign hdmi_out0_dram_port_cmd_fifo_asyncfifo_dout = hdmi_out0_dram_port_cmd_fifo_rdport_dat_r;
always @(*) begin
	hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary <= 3'd0;
	if (hdmi_out0_dram_port_cmd_fifo_graycounter0_ce) begin
		hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary <= (hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary <= hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary;
	end
end
assign hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next = (hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary ^ hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary[2:1]);
always @(*) begin
	hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary <= 3'd0;
	if (hdmi_out0_dram_port_cmd_fifo_graycounter1_ce) begin
		hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary <= (hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary <= hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary;
	end
end
assign hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next = (hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary ^ hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary[2:1]);
assign hdmi_out0_dram_port_cmd_fifo_sink_valid = hdmi_out0_dram_port_litedramport0_cmd_valid;
assign hdmi_out0_dram_port_litedramport0_cmd_ready = hdmi_out0_dram_port_cmd_fifo_sink_ready;
assign hdmi_out0_dram_port_cmd_fifo_sink_first = hdmi_out0_dram_port_litedramport0_cmd_first;
assign hdmi_out0_dram_port_cmd_fifo_sink_last = hdmi_out0_dram_port_litedramport0_cmd_last;
assign hdmi_out0_dram_port_cmd_fifo_sink_payload_we = hdmi_out0_dram_port_litedramport0_cmd_payload_we;
assign hdmi_out0_dram_port_cmd_fifo_sink_payload_adr = hdmi_out0_dram_port_litedramport0_cmd_payload_adr;
assign hdmi_out0_dram_port_cmd_valid = hdmi_out0_dram_port_cmd_fifo_source_valid;
assign hdmi_out0_dram_port_cmd_fifo_source_ready = hdmi_out0_dram_port_cmd_ready;
assign hdmi_out0_dram_port_cmd_first = hdmi_out0_dram_port_cmd_fifo_source_first;
assign hdmi_out0_dram_port_cmd_last = hdmi_out0_dram_port_cmd_fifo_source_last;
assign hdmi_out0_dram_port_cmd_payload_we = hdmi_out0_dram_port_cmd_fifo_source_payload_we;
assign hdmi_out0_dram_port_cmd_payload_adr = hdmi_out0_dram_port_cmd_fifo_source_payload_adr;
assign hdmi_out0_dram_port_rdata_fifo_asyncfifo_din = {hdmi_out0_dram_port_rdata_fifo_fifo_in_last, hdmi_out0_dram_port_rdata_fifo_fifo_in_first, hdmi_out0_dram_port_rdata_fifo_fifo_in_payload_data};
assign {hdmi_out0_dram_port_rdata_fifo_fifo_out_last, hdmi_out0_dram_port_rdata_fifo_fifo_out_first, hdmi_out0_dram_port_rdata_fifo_fifo_out_payload_data} = hdmi_out0_dram_port_rdata_fifo_asyncfifo_dout;
assign hdmi_out0_dram_port_rdata_fifo_sink_ready = hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable;
assign hdmi_out0_dram_port_rdata_fifo_asyncfifo_we = hdmi_out0_dram_port_rdata_fifo_sink_valid;
assign hdmi_out0_dram_port_rdata_fifo_fifo_in_first = hdmi_out0_dram_port_rdata_fifo_sink_first;
assign hdmi_out0_dram_port_rdata_fifo_fifo_in_last = hdmi_out0_dram_port_rdata_fifo_sink_last;
assign hdmi_out0_dram_port_rdata_fifo_fifo_in_payload_data = hdmi_out0_dram_port_rdata_fifo_sink_payload_data;
assign hdmi_out0_dram_port_rdata_fifo_source_valid = hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable;
assign hdmi_out0_dram_port_rdata_fifo_source_first = hdmi_out0_dram_port_rdata_fifo_fifo_out_first;
assign hdmi_out0_dram_port_rdata_fifo_source_last = hdmi_out0_dram_port_rdata_fifo_fifo_out_last;
assign hdmi_out0_dram_port_rdata_fifo_source_payload_data = hdmi_out0_dram_port_rdata_fifo_fifo_out_payload_data;
assign hdmi_out0_dram_port_rdata_fifo_asyncfifo_re = hdmi_out0_dram_port_rdata_fifo_source_ready;
assign hdmi_out0_dram_port_rdata_fifo_graycounter0_ce = (hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable & hdmi_out0_dram_port_rdata_fifo_asyncfifo_we);
assign hdmi_out0_dram_port_rdata_fifo_graycounter1_ce = (hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable & hdmi_out0_dram_port_rdata_fifo_asyncfifo_re);
assign hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable = (((hdmi_out0_dram_port_rdata_fifo_graycounter0_q[4] == hdmi_out0_dram_port_rdata_fifo_consume_wdomain[4]) | (hdmi_out0_dram_port_rdata_fifo_graycounter0_q[3] == hdmi_out0_dram_port_rdata_fifo_consume_wdomain[3])) | (hdmi_out0_dram_port_rdata_fifo_graycounter0_q[2:0] != hdmi_out0_dram_port_rdata_fifo_consume_wdomain[2:0]));
assign hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable = (hdmi_out0_dram_port_rdata_fifo_graycounter1_q != hdmi_out0_dram_port_rdata_fifo_produce_rdomain);
assign hdmi_out0_dram_port_rdata_fifo_wrport_adr = hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary[3:0];
assign hdmi_out0_dram_port_rdata_fifo_wrport_dat_w = hdmi_out0_dram_port_rdata_fifo_asyncfifo_din;
assign hdmi_out0_dram_port_rdata_fifo_wrport_we = hdmi_out0_dram_port_rdata_fifo_graycounter0_ce;
assign hdmi_out0_dram_port_rdata_fifo_rdport_adr = hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary[3:0];
assign hdmi_out0_dram_port_rdata_fifo_asyncfifo_dout = hdmi_out0_dram_port_rdata_fifo_rdport_dat_r;
always @(*) begin
	hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary <= 5'd0;
	if (hdmi_out0_dram_port_rdata_fifo_graycounter0_ce) begin
		hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary <= (hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary <= hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary;
	end
end
assign hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next = (hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary ^ hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary[4:1]);
always @(*) begin
	hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary <= 5'd0;
	if (hdmi_out0_dram_port_rdata_fifo_graycounter1_ce) begin
		hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary <= (hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary <= hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary;
	end
end
assign hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next = (hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary ^ hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary[4:1]);
assign hdmi_out0_dram_port_rdata_fifo_sink_valid = hdmi_out0_dram_port_rdata_valid;
assign hdmi_out0_dram_port_rdata_ready = hdmi_out0_dram_port_rdata_fifo_sink_ready;
assign hdmi_out0_dram_port_rdata_fifo_sink_first = hdmi_out0_dram_port_rdata_first;
assign hdmi_out0_dram_port_rdata_fifo_sink_last = hdmi_out0_dram_port_rdata_last;
assign hdmi_out0_dram_port_rdata_fifo_sink_payload_data = hdmi_out0_dram_port_rdata_payload_data;
assign hdmi_out0_dram_port_litedramport0_rdata_valid = hdmi_out0_dram_port_rdata_fifo_source_valid;
assign hdmi_out0_dram_port_rdata_fifo_source_ready = hdmi_out0_dram_port_litedramport0_rdata_ready;
assign hdmi_out0_dram_port_litedramport0_rdata_first = hdmi_out0_dram_port_rdata_fifo_source_first;
assign hdmi_out0_dram_port_litedramport0_rdata_last = hdmi_out0_dram_port_rdata_fifo_source_last;
assign hdmi_out0_dram_port_litedramport0_rdata_payload_data = hdmi_out0_dram_port_rdata_fifo_source_payload_data;
always @(*) begin
	hdmi_out0_dram_port_litedramport1_cmd_ready <= 1'd0;
	hdmi_out0_dram_port_counter_ce <= 1'd0;
	hdmi_out0_dram_port_litedramport0_cmd_valid <= 1'd0;
	hdmi_out0_dram_port_litedramport0_cmd_payload_adr <= 25'd0;
	if (hdmi_out0_dram_port_litedramport1_cmd_valid) begin
		if ((hdmi_out0_dram_port_counter == 1'd0)) begin
			hdmi_out0_dram_port_litedramport0_cmd_valid <= 1'd1;
			hdmi_out0_dram_port_litedramport0_cmd_payload_adr <= hdmi_out0_dram_port_litedramport1_cmd_payload_adr[27:3];
			hdmi_out0_dram_port_litedramport1_cmd_ready <= hdmi_out0_dram_port_litedramport0_cmd_ready;
			hdmi_out0_dram_port_counter_ce <= hdmi_out0_dram_port_litedramport0_cmd_ready;
		end else begin
			hdmi_out0_dram_port_litedramport1_cmd_ready <= 1'd1;
			hdmi_out0_dram_port_counter_ce <= 1'd1;
		end
	end
end
always @(*) begin
	hdmi_out0_dram_port_cmd_buffer_sink_valid <= 1'd0;
	hdmi_out0_dram_port_cmd_buffer_sink_payload_sel <= 8'd0;
	if ((hdmi_out0_dram_port_litedramport0_cmd_valid & hdmi_out0_dram_port_litedramport0_cmd_ready)) begin
		hdmi_out0_dram_port_cmd_buffer_sink_valid <= 1'd1;
		hdmi_out0_dram_port_cmd_buffer_sink_payload_sel <= 8'd255;
	end
end
assign hdmi_out0_dram_port_rdata_buffer_sink_valid = hdmi_out0_dram_port_litedramport0_rdata_valid;
assign hdmi_out0_dram_port_litedramport0_rdata_ready = hdmi_out0_dram_port_rdata_buffer_sink_ready;
assign hdmi_out0_dram_port_rdata_buffer_sink_first = hdmi_out0_dram_port_litedramport0_rdata_first;
assign hdmi_out0_dram_port_rdata_buffer_sink_last = hdmi_out0_dram_port_litedramport0_rdata_last;
assign hdmi_out0_dram_port_rdata_buffer_sink_payload_data = hdmi_out0_dram_port_litedramport0_rdata_payload_data;
assign hdmi_out0_dram_port_rdata_converter_sink_valid = hdmi_out0_dram_port_rdata_buffer_source_valid;
assign hdmi_out0_dram_port_rdata_buffer_source_ready = hdmi_out0_dram_port_rdata_converter_sink_ready;
assign hdmi_out0_dram_port_rdata_converter_sink_first = hdmi_out0_dram_port_rdata_buffer_source_first;
assign hdmi_out0_dram_port_rdata_converter_sink_last = hdmi_out0_dram_port_rdata_buffer_source_last;
assign hdmi_out0_dram_port_rdata_converter_sink_payload_data = hdmi_out0_dram_port_rdata_buffer_source_payload_data;
assign hdmi_out0_dram_port_rdata_chunk_valid = ((hdmi_out0_dram_port_cmd_buffer_source_payload_sel & hdmi_out0_dram_port_rdata_chunk) != 1'd0);
always @(*) begin
	hdmi_out0_dram_port_rdata_converter_source_ready <= 1'd0;
	hdmi_out0_dram_port_litedramport1_rdata_payload_data <= 16'd0;
	hdmi_out0_dram_port_litedramport1_rdata_valid <= 1'd0;
	if (hdmi_out0_dram_port_litedramport1_flush) begin
		hdmi_out0_dram_port_rdata_converter_source_ready <= 1'd1;
	end else begin
		if (hdmi_out0_dram_port_cmd_buffer_source_valid) begin
			if (hdmi_out0_dram_port_rdata_chunk_valid) begin
				hdmi_out0_dram_port_litedramport1_rdata_valid <= hdmi_out0_dram_port_rdata_converter_source_valid;
				hdmi_out0_dram_port_litedramport1_rdata_payload_data <= hdmi_out0_dram_port_rdata_converter_source_payload_data;
				hdmi_out0_dram_port_rdata_converter_source_ready <= hdmi_out0_dram_port_litedramport1_rdata_ready;
			end else begin
				hdmi_out0_dram_port_rdata_converter_source_ready <= 1'd1;
			end
		end
	end
end
assign hdmi_out0_dram_port_cmd_buffer_source_ready = (hdmi_out0_dram_port_rdata_converter_source_ready & hdmi_out0_dram_port_rdata_chunk[7]);
assign hdmi_out0_dram_port_cmd_buffer_syncfifo_din = {hdmi_out0_dram_port_cmd_buffer_fifo_in_last, hdmi_out0_dram_port_cmd_buffer_fifo_in_first, hdmi_out0_dram_port_cmd_buffer_fifo_in_payload_sel};
assign {hdmi_out0_dram_port_cmd_buffer_fifo_out_last, hdmi_out0_dram_port_cmd_buffer_fifo_out_first, hdmi_out0_dram_port_cmd_buffer_fifo_out_payload_sel} = hdmi_out0_dram_port_cmd_buffer_syncfifo_dout;
assign hdmi_out0_dram_port_cmd_buffer_sink_ready = hdmi_out0_dram_port_cmd_buffer_syncfifo_writable;
assign hdmi_out0_dram_port_cmd_buffer_syncfifo_we = hdmi_out0_dram_port_cmd_buffer_sink_valid;
assign hdmi_out0_dram_port_cmd_buffer_fifo_in_first = hdmi_out0_dram_port_cmd_buffer_sink_first;
assign hdmi_out0_dram_port_cmd_buffer_fifo_in_last = hdmi_out0_dram_port_cmd_buffer_sink_last;
assign hdmi_out0_dram_port_cmd_buffer_fifo_in_payload_sel = hdmi_out0_dram_port_cmd_buffer_sink_payload_sel;
assign hdmi_out0_dram_port_cmd_buffer_source_valid = hdmi_out0_dram_port_cmd_buffer_syncfifo_readable;
assign hdmi_out0_dram_port_cmd_buffer_source_first = hdmi_out0_dram_port_cmd_buffer_fifo_out_first;
assign hdmi_out0_dram_port_cmd_buffer_source_last = hdmi_out0_dram_port_cmd_buffer_fifo_out_last;
assign hdmi_out0_dram_port_cmd_buffer_source_payload_sel = hdmi_out0_dram_port_cmd_buffer_fifo_out_payload_sel;
assign hdmi_out0_dram_port_cmd_buffer_syncfifo_re = hdmi_out0_dram_port_cmd_buffer_source_ready;
always @(*) begin
	hdmi_out0_dram_port_cmd_buffer_wrport_adr <= 2'd0;
	if (hdmi_out0_dram_port_cmd_buffer_replace) begin
		hdmi_out0_dram_port_cmd_buffer_wrport_adr <= (hdmi_out0_dram_port_cmd_buffer_produce - 1'd1);
	end else begin
		hdmi_out0_dram_port_cmd_buffer_wrport_adr <= hdmi_out0_dram_port_cmd_buffer_produce;
	end
end
assign hdmi_out0_dram_port_cmd_buffer_wrport_dat_w = hdmi_out0_dram_port_cmd_buffer_syncfifo_din;
assign hdmi_out0_dram_port_cmd_buffer_wrport_we = (hdmi_out0_dram_port_cmd_buffer_syncfifo_we & (hdmi_out0_dram_port_cmd_buffer_syncfifo_writable | hdmi_out0_dram_port_cmd_buffer_replace));
assign hdmi_out0_dram_port_cmd_buffer_do_read = (hdmi_out0_dram_port_cmd_buffer_syncfifo_readable & hdmi_out0_dram_port_cmd_buffer_syncfifo_re);
assign hdmi_out0_dram_port_cmd_buffer_rdport_adr = hdmi_out0_dram_port_cmd_buffer_consume;
assign hdmi_out0_dram_port_cmd_buffer_syncfifo_dout = hdmi_out0_dram_port_cmd_buffer_rdport_dat_r;
assign hdmi_out0_dram_port_cmd_buffer_syncfifo_writable = (hdmi_out0_dram_port_cmd_buffer_level != 3'd4);
assign hdmi_out0_dram_port_cmd_buffer_syncfifo_readable = (hdmi_out0_dram_port_cmd_buffer_level != 1'd0);
assign hdmi_out0_dram_port_rdata_buffer_pipe_ce = (hdmi_out0_dram_port_rdata_buffer_source_ready | (~hdmi_out0_dram_port_rdata_buffer_valid_n));
assign hdmi_out0_dram_port_rdata_buffer_sink_ready = hdmi_out0_dram_port_rdata_buffer_pipe_ce;
assign hdmi_out0_dram_port_rdata_buffer_source_valid = hdmi_out0_dram_port_rdata_buffer_valid_n;
assign hdmi_out0_dram_port_rdata_buffer_busy = (1'd0 | hdmi_out0_dram_port_rdata_buffer_valid_n);
assign hdmi_out0_dram_port_rdata_buffer_source_first = hdmi_out0_dram_port_rdata_buffer_first_n;
assign hdmi_out0_dram_port_rdata_buffer_source_last = hdmi_out0_dram_port_rdata_buffer_last_n;
assign hdmi_out0_dram_port_rdata_converter_converter_sink_valid = hdmi_out0_dram_port_rdata_converter_sink_valid;
assign hdmi_out0_dram_port_rdata_converter_converter_sink_first = hdmi_out0_dram_port_rdata_converter_sink_first;
assign hdmi_out0_dram_port_rdata_converter_converter_sink_last = hdmi_out0_dram_port_rdata_converter_sink_last;
assign hdmi_out0_dram_port_rdata_converter_sink_ready = hdmi_out0_dram_port_rdata_converter_converter_sink_ready;
always @(*) begin
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data <= 128'd0;
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[15:0] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[15:0];
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[31:16] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[31:16];
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[47:32] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[47:32];
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[63:48] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[63:48];
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[79:64] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[79:64];
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[95:80] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[95:80];
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[111:96] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[111:96];
	hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[127:112] <= hdmi_out0_dram_port_rdata_converter_sink_payload_data[127:112];
end
assign hdmi_out0_dram_port_rdata_converter_source_valid = hdmi_out0_dram_port_rdata_converter_source_source_valid;
assign hdmi_out0_dram_port_rdata_converter_source_first = hdmi_out0_dram_port_rdata_converter_source_source_first;
assign hdmi_out0_dram_port_rdata_converter_source_last = hdmi_out0_dram_port_rdata_converter_source_source_last;
assign hdmi_out0_dram_port_rdata_converter_source_source_ready = hdmi_out0_dram_port_rdata_converter_source_ready;
assign {hdmi_out0_dram_port_rdata_converter_source_payload_data} = hdmi_out0_dram_port_rdata_converter_source_source_payload_data;
assign hdmi_out0_dram_port_rdata_converter_source_source_valid = hdmi_out0_dram_port_rdata_converter_converter_source_valid;
assign hdmi_out0_dram_port_rdata_converter_converter_source_ready = hdmi_out0_dram_port_rdata_converter_source_source_ready;
assign hdmi_out0_dram_port_rdata_converter_source_source_first = hdmi_out0_dram_port_rdata_converter_converter_source_first;
assign hdmi_out0_dram_port_rdata_converter_source_source_last = hdmi_out0_dram_port_rdata_converter_converter_source_last;
assign hdmi_out0_dram_port_rdata_converter_source_source_payload_data = hdmi_out0_dram_port_rdata_converter_converter_source_payload_data;
assign hdmi_out0_dram_port_rdata_converter_converter_first = (hdmi_out0_dram_port_rdata_converter_converter_mux == 1'd0);
assign hdmi_out0_dram_port_rdata_converter_converter_last = (hdmi_out0_dram_port_rdata_converter_converter_mux == 3'd7);
assign hdmi_out0_dram_port_rdata_converter_converter_source_valid = hdmi_out0_dram_port_rdata_converter_converter_sink_valid;
assign hdmi_out0_dram_port_rdata_converter_converter_source_first = (hdmi_out0_dram_port_rdata_converter_converter_sink_first & hdmi_out0_dram_port_rdata_converter_converter_first);
assign hdmi_out0_dram_port_rdata_converter_converter_source_last = (hdmi_out0_dram_port_rdata_converter_converter_sink_last & hdmi_out0_dram_port_rdata_converter_converter_last);
assign hdmi_out0_dram_port_rdata_converter_converter_sink_ready = (hdmi_out0_dram_port_rdata_converter_converter_last & hdmi_out0_dram_port_rdata_converter_converter_source_ready);
always @(*) begin
	hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= 16'd0;
	case (hdmi_out0_dram_port_rdata_converter_converter_mux)
		1'd0: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[127:112];
		end
		1'd1: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[111:96];
		end
		2'd2: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[95:80];
		end
		2'd3: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[79:64];
		end
		3'd4: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[63:48];
		end
		3'd5: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[47:32];
		end
		3'd6: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[31:16];
		end
		default: begin
			hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[15:0];
		end
	endcase
end
assign hdmi_out0_dram_port_rdata_converter_converter_source_payload_valid_token_count = hdmi_out0_dram_port_rdata_converter_converter_last;
assign videosoc_data_port_adr = videosoc_interface0_wb_sdram_adr[10:2];
always @(*) begin
	videosoc_data_port_dat_w <= 128'd0;
	videosoc_data_port_we <= 16'd0;
	if (videosoc_write_from_slave) begin
		videosoc_data_port_dat_w <= videosoc_interface_dat_r;
		videosoc_data_port_we <= {16{1'd1}};
	end else begin
		videosoc_data_port_dat_w <= {4{videosoc_interface0_wb_sdram_dat_w}};
		if ((((videosoc_interface0_wb_sdram_cyc & videosoc_interface0_wb_sdram_stb) & videosoc_interface0_wb_sdram_we) & videosoc_interface0_wb_sdram_ack)) begin
			videosoc_data_port_we <= {({4{(videosoc_interface0_wb_sdram_adr[1:0] == 1'd0)}} & videosoc_interface0_wb_sdram_sel), ({4{(videosoc_interface0_wb_sdram_adr[1:0] == 1'd1)}} & videosoc_interface0_wb_sdram_sel), ({4{(videosoc_interface0_wb_sdram_adr[1:0] == 2'd2)}} & videosoc_interface0_wb_sdram_sel), ({4{(videosoc_interface0_wb_sdram_adr[1:0] == 2'd3)}} & videosoc_interface0_wb_sdram_sel)};
		end
	end
end
assign videosoc_interface_dat_w = videosoc_data_port_dat_r;
assign videosoc_interface_sel = 16'd65535;
always @(*) begin
	videosoc_interface0_wb_sdram_dat_r <= 32'd0;
	case (videosoc_adr_offset_r)
		1'd0: begin
			videosoc_interface0_wb_sdram_dat_r <= videosoc_data_port_dat_r[127:96];
		end
		1'd1: begin
			videosoc_interface0_wb_sdram_dat_r <= videosoc_data_port_dat_r[95:64];
		end
		2'd2: begin
			videosoc_interface0_wb_sdram_dat_r <= videosoc_data_port_dat_r[63:32];
		end
		default: begin
			videosoc_interface0_wb_sdram_dat_r <= videosoc_data_port_dat_r[31:0];
		end
	endcase
end
assign {videosoc_tag_do_dirty, videosoc_tag_do_tag} = videosoc_tag_port_dat_r;
assign videosoc_tag_port_dat_w = {videosoc_tag_di_dirty, videosoc_tag_di_tag};
assign videosoc_tag_port_adr = videosoc_interface0_wb_sdram_adr[10:2];
assign videosoc_tag_di_tag = videosoc_interface0_wb_sdram_adr[29:11];
assign videosoc_interface_adr = {videosoc_tag_do_tag, videosoc_interface0_wb_sdram_adr[10:2]};
always @(*) begin
	videosoc_word_inc <= 1'd0;
	videosoc_write_from_slave <= 1'd0;
	videosoc_interface_cyc <= 1'd0;
	videosoc_interface_stb <= 1'd0;
	videosoc_tag_port_we <= 1'd0;
	videosoc_interface0_wb_sdram_ack <= 1'd0;
	videosoc_interface_we <= 1'd0;
	fullmemorywe_next_state <= 3'd0;
	videosoc_tag_di_dirty <= 1'd0;
	videosoc_word_clr <= 1'd0;
	fullmemorywe_next_state <= fullmemorywe_state;
	case (fullmemorywe_state)
		1'd1: begin
			videosoc_word_clr <= 1'd1;
			if ((videosoc_tag_do_tag == videosoc_interface0_wb_sdram_adr[29:11])) begin
				videosoc_interface0_wb_sdram_ack <= 1'd1;
				if (videosoc_interface0_wb_sdram_we) begin
					videosoc_tag_di_dirty <= 1'd1;
					videosoc_tag_port_we <= 1'd1;
				end
				fullmemorywe_next_state <= 1'd0;
			end else begin
				if (videosoc_tag_do_dirty) begin
					fullmemorywe_next_state <= 2'd2;
				end else begin
					fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			videosoc_interface_stb <= 1'd1;
			videosoc_interface_cyc <= 1'd1;
			videosoc_interface_we <= 1'd1;
			if (videosoc_interface_ack) begin
				videosoc_word_inc <= 1'd1;
				if (1'd1) begin
					fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			videosoc_tag_port_we <= 1'd1;
			videosoc_word_clr <= 1'd1;
			fullmemorywe_next_state <= 3'd4;
		end
		3'd4: begin
			videosoc_interface_stb <= 1'd1;
			videosoc_interface_cyc <= 1'd1;
			videosoc_interface_we <= 1'd0;
			if (videosoc_interface_ack) begin
				videosoc_write_from_slave <= 1'd1;
				videosoc_word_inc <= 1'd1;
				if (1'd1) begin
					fullmemorywe_next_state <= 1'd1;
				end else begin
					fullmemorywe_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((videosoc_interface0_wb_sdram_cyc & videosoc_interface0_wb_sdram_stb)) begin
				fullmemorywe_next_state <= 1'd1;
			end
		end
	endcase
end
assign videosoc_port_cmd_payload_adr = videosoc_interface_adr;
assign videosoc_port_wdata_payload_we = videosoc_interface_sel;
assign videosoc_port_wdata_payload_data = videosoc_interface_dat_w;
assign videosoc_interface_dat_r = videosoc_port_rdata_payload_data;
always @(*) begin
	videosoc_port_cmd_valid <= 1'd0;
	videosoc_port_cmd_payload_we <= 1'd0;
	videosoc_port_rdata_ready <= 1'd0;
	videosoc_port_wdata_valid <= 1'd0;
	litedramwishbonebridge_next_state <= 2'd0;
	videosoc_interface_ack <= 1'd0;
	litedramwishbonebridge_next_state <= litedramwishbonebridge_state;
	case (litedramwishbonebridge_state)
		1'd1: begin
			videosoc_port_cmd_valid <= 1'd1;
			videosoc_port_cmd_payload_we <= videosoc_interface_we;
			if (videosoc_port_cmd_ready) begin
				if (videosoc_interface_we) begin
					litedramwishbonebridge_next_state <= 2'd2;
				end else begin
					litedramwishbonebridge_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			videosoc_port_wdata_valid <= 1'd1;
			if (videosoc_port_wdata_ready) begin
				videosoc_interface_ack <= 1'd1;
				litedramwishbonebridge_next_state <= 1'd0;
			end
		end
		2'd3: begin
			videosoc_port_rdata_ready <= 1'd1;
			if (videosoc_port_rdata_valid) begin
				videosoc_interface_ack <= 1'd1;
				litedramwishbonebridge_next_state <= 1'd0;
			end
		end
		default: begin
			if ((videosoc_interface_cyc & videosoc_interface_stb)) begin
				litedramwishbonebridge_next_state <= 1'd1;
			end
		end
	endcase
end
assign spiflash_1x_wp = 1'd1;
assign spiflash_1x_hold = 1'd1;
assign videosoc_bus_dat_r = videosoc_sr;
always @(*) begin
	videosoc_miso_status <= 1'd0;
	spiflash_1x_mosi <= 1'd0;
	spiflash_1x_cs_n <= 1'd0;
	videosoc_clk0 <= 1'd0;
	if (videosoc_bitbang_en_storage) begin
		videosoc_clk0 <= videosoc_bitbang_storage[1];
		spiflash_1x_cs_n <= videosoc_bitbang_storage[2];
		if (videosoc_bitbang_storage[1]) begin
			videosoc_miso_status <= spiflash_1x_miso;
		end
		spiflash_1x_mosi <= videosoc_bitbang_storage[0];
	end else begin
		videosoc_clk0 <= videosoc_clk1;
		spiflash_1x_cs_n <= videosoc_cs_n;
		spiflash_1x_mosi <= videosoc_sr[31];
	end
end
assign ethphy_reset0 = (ethphy_reset_storage | ethphy_reset1);
assign eth_rst_n = (~ethphy_reset0);
assign ethphy_counter_done = (ethphy_counter == 9'd256);
assign ethphy_counter_ce = (~ethphy_counter_done);
assign ethphy_reset1 = (~ethphy_counter_done);
assign ethphy_sink_ready = 1'd1;
assign ethphy_last = ((~ethphy_rx_ctl) & ethphy_rx_ctl_d);
assign ethphy_source_last = ethphy_last;
assign eth_mdc = ethphy_storage[0];
assign ethphy_data_oe = ethphy_storage[1];
assign ethphy_data_w = ethphy_storage[2];
assign ethmac_tx_cdc_sink_valid = ethmac_source_valid;
assign ethmac_source_ready = ethmac_tx_cdc_sink_ready;
assign ethmac_tx_cdc_sink_first = ethmac_source_first;
assign ethmac_tx_cdc_sink_last = ethmac_source_last;
assign ethmac_tx_cdc_sink_payload_data = ethmac_source_payload_data;
assign ethmac_tx_cdc_sink_payload_last_be = ethmac_source_payload_last_be;
assign ethmac_tx_cdc_sink_payload_error = ethmac_source_payload_error;
assign ethmac_sink_valid = ethmac_rx_cdc_source_valid;
assign ethmac_rx_cdc_source_ready = ethmac_sink_ready;
assign ethmac_sink_first = ethmac_rx_cdc_source_first;
assign ethmac_sink_last = ethmac_rx_cdc_source_last;
assign ethmac_sink_payload_data = ethmac_rx_cdc_source_payload_data;
assign ethmac_sink_payload_last_be = ethmac_rx_cdc_source_payload_last_be;
assign ethmac_sink_payload_error = ethmac_rx_cdc_source_payload_error;
assign ethmac_ps_preamble_error_i = ethmac_preamble_checker_error;
assign ethmac_ps_crc_error_i = ethmac_crc32_checker_error;
always @(*) begin
	ethmac_tx_gap_inserter_source_payload_error <= 1'd0;
	ethmac_tx_gap_inserter_counter_reset <= 1'd0;
	ethmac_tx_gap_inserter_source_payload_data <= 8'd0;
	ethmac_tx_gap_inserter_counter_ce <= 1'd0;
	ethmac_tx_gap_inserter_sink_ready <= 1'd0;
	ethmac_tx_gap_inserter_source_valid <= 1'd0;
	ethmac_tx_gap_inserter_source_first <= 1'd0;
	ethmac_tx_gap_inserter_source_last <= 1'd0;
	liteethmacgap_next_state <= 1'd0;
	ethmac_tx_gap_inserter_source_payload_last_be <= 1'd0;
	liteethmacgap_next_state <= liteethmacgap_state;
	case (liteethmacgap_state)
		1'd1: begin
			ethmac_tx_gap_inserter_counter_ce <= 1'd1;
			if ((ethmac_tx_gap_inserter_counter == 4'd11)) begin
				liteethmacgap_next_state <= 1'd0;
			end
		end
		default: begin
			ethmac_tx_gap_inserter_counter_reset <= 1'd1;
			ethmac_tx_gap_inserter_source_valid <= ethmac_tx_gap_inserter_sink_valid;
			ethmac_tx_gap_inserter_sink_ready <= ethmac_tx_gap_inserter_source_ready;
			ethmac_tx_gap_inserter_source_first <= ethmac_tx_gap_inserter_sink_first;
			ethmac_tx_gap_inserter_source_last <= ethmac_tx_gap_inserter_sink_last;
			ethmac_tx_gap_inserter_source_payload_data <= ethmac_tx_gap_inserter_sink_payload_data;
			ethmac_tx_gap_inserter_source_payload_last_be <= ethmac_tx_gap_inserter_sink_payload_last_be;
			ethmac_tx_gap_inserter_source_payload_error <= ethmac_tx_gap_inserter_sink_payload_error;
			if (((ethmac_tx_gap_inserter_sink_valid & ethmac_tx_gap_inserter_sink_last) & ethmac_tx_gap_inserter_sink_ready)) begin
				liteethmacgap_next_state <= 1'd1;
			end
		end
	endcase
end
assign ethmac_preamble_inserter_source_payload_last_be = ethmac_preamble_inserter_sink_payload_last_be;
always @(*) begin
	ethmac_preamble_inserter_inc_cnt <= 1'd0;
	ethmac_preamble_inserter_source_valid <= 1'd0;
	liteethmacpreambleinserter_next_state <= 2'd0;
	ethmac_preamble_inserter_source_first <= 1'd0;
	ethmac_preamble_inserter_source_last <= 1'd0;
	ethmac_preamble_inserter_source_payload_data <= 8'd0;
	ethmac_preamble_inserter_source_payload_error <= 1'd0;
	ethmac_preamble_inserter_clr_cnt <= 1'd0;
	ethmac_preamble_inserter_sink_ready <= 1'd0;
	ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_sink_payload_data;
	liteethmacpreambleinserter_next_state <= liteethmacpreambleinserter_state;
	case (liteethmacpreambleinserter_state)
		1'd1: begin
			ethmac_preamble_inserter_source_valid <= 1'd1;
			case (ethmac_preamble_inserter_cnt)
				1'd0: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[7:0];
				end
				1'd1: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[15:8];
				end
				2'd2: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[23:16];
				end
				2'd3: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[31:24];
				end
				3'd4: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[39:32];
				end
				3'd5: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[47:40];
				end
				3'd6: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[55:48];
				end
				default: begin
					ethmac_preamble_inserter_source_payload_data <= ethmac_preamble_inserter_preamble[63:56];
				end
			endcase
			if ((ethmac_preamble_inserter_cnt == 3'd7)) begin
				if (ethmac_preamble_inserter_source_ready) begin
					liteethmacpreambleinserter_next_state <= 2'd2;
				end
			end else begin
				ethmac_preamble_inserter_inc_cnt <= ethmac_preamble_inserter_source_ready;
			end
		end
		2'd2: begin
			ethmac_preamble_inserter_source_valid <= ethmac_preamble_inserter_sink_valid;
			ethmac_preamble_inserter_sink_ready <= ethmac_preamble_inserter_source_ready;
			ethmac_preamble_inserter_source_first <= ethmac_preamble_inserter_sink_first;
			ethmac_preamble_inserter_source_last <= ethmac_preamble_inserter_sink_last;
			ethmac_preamble_inserter_source_payload_error <= ethmac_preamble_inserter_sink_payload_error;
			if (((ethmac_preamble_inserter_sink_valid & ethmac_preamble_inserter_sink_last) & ethmac_preamble_inserter_source_ready)) begin
				liteethmacpreambleinserter_next_state <= 1'd0;
			end
		end
		default: begin
			ethmac_preamble_inserter_sink_ready <= 1'd1;
			ethmac_preamble_inserter_clr_cnt <= 1'd1;
			if (ethmac_preamble_inserter_sink_valid) begin
				ethmac_preamble_inserter_sink_ready <= 1'd0;
				liteethmacpreambleinserter_next_state <= 1'd1;
			end
		end
	endcase
end
assign ethmac_preamble_checker_source_payload_data = ethmac_preamble_checker_sink_payload_data;
assign ethmac_preamble_checker_source_payload_last_be = ethmac_preamble_checker_sink_payload_last_be;
always @(*) begin
	liteethmacpreamblechecker_next_state <= 1'd0;
	ethmac_preamble_checker_source_payload_error <= 1'd0;
	ethmac_preamble_checker_sink_ready <= 1'd0;
	ethmac_preamble_checker_error <= 1'd0;
	ethmac_preamble_checker_source_valid <= 1'd0;
	ethmac_preamble_checker_source_first <= 1'd0;
	ethmac_preamble_checker_source_last <= 1'd0;
	liteethmacpreamblechecker_next_state <= liteethmacpreamblechecker_state;
	case (liteethmacpreamblechecker_state)
		1'd1: begin
			ethmac_preamble_checker_source_valid <= ethmac_preamble_checker_sink_valid;
			ethmac_preamble_checker_sink_ready <= ethmac_preamble_checker_source_ready;
			ethmac_preamble_checker_source_first <= ethmac_preamble_checker_sink_first;
			ethmac_preamble_checker_source_last <= ethmac_preamble_checker_sink_last;
			ethmac_preamble_checker_source_payload_error <= ethmac_preamble_checker_sink_payload_error;
			if (((ethmac_preamble_checker_source_valid & ethmac_preamble_checker_source_last) & ethmac_preamble_checker_source_ready)) begin
				liteethmacpreamblechecker_next_state <= 1'd0;
			end
		end
		default: begin
			ethmac_preamble_checker_sink_ready <= 1'd1;
			if (((ethmac_preamble_checker_sink_valid & (~ethmac_preamble_checker_sink_last)) & (ethmac_preamble_checker_sink_payload_data == 8'd213))) begin
				liteethmacpreamblechecker_next_state <= 1'd1;
			end
			if ((ethmac_preamble_checker_sink_valid & ethmac_preamble_checker_sink_last)) begin
				ethmac_preamble_checker_error <= 1'd1;
			end
		end
	endcase
end
assign ethmac_crc32_inserter_cnt_done = (ethmac_crc32_inserter_cnt == 1'd0);
assign ethmac_crc32_inserter_data1 = ethmac_crc32_inserter_data0;
assign ethmac_crc32_inserter_last = ethmac_crc32_inserter_reg;
assign ethmac_crc32_inserter_value = (~{ethmac_crc32_inserter_reg[0], ethmac_crc32_inserter_reg[1], ethmac_crc32_inserter_reg[2], ethmac_crc32_inserter_reg[3], ethmac_crc32_inserter_reg[4], ethmac_crc32_inserter_reg[5], ethmac_crc32_inserter_reg[6], ethmac_crc32_inserter_reg[7], ethmac_crc32_inserter_reg[8], ethmac_crc32_inserter_reg[9], ethmac_crc32_inserter_reg[10], ethmac_crc32_inserter_reg[11], ethmac_crc32_inserter_reg[12], ethmac_crc32_inserter_reg[13], ethmac_crc32_inserter_reg[14], ethmac_crc32_inserter_reg[15], ethmac_crc32_inserter_reg[16], ethmac_crc32_inserter_reg[17], ethmac_crc32_inserter_reg[18], ethmac_crc32_inserter_reg[19], ethmac_crc32_inserter_reg[20], ethmac_crc32_inserter_reg[21], ethmac_crc32_inserter_reg[22], ethmac_crc32_inserter_reg[23], ethmac_crc32_inserter_reg[24], ethmac_crc32_inserter_reg[25], ethmac_crc32_inserter_reg[26], ethmac_crc32_inserter_reg[27], ethmac_crc32_inserter_reg[28], ethmac_crc32_inserter_reg[29], ethmac_crc32_inserter_reg[30], ethmac_crc32_inserter_reg[31]});
assign ethmac_crc32_inserter_error = (ethmac_crc32_inserter_next != 32'd3338984827);
always @(*) begin
	ethmac_crc32_inserter_next <= 32'd0;
	ethmac_crc32_inserter_next[0] <= (((ethmac_crc32_inserter_last[24] ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[1] <= (((((((ethmac_crc32_inserter_last[25] ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[2] <= (((((((((ethmac_crc32_inserter_last[26] ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[3] <= (((((((ethmac_crc32_inserter_last[27] ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]);
	ethmac_crc32_inserter_next[4] <= (((((((((ethmac_crc32_inserter_last[28] ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[5] <= (((((((((((((ethmac_crc32_inserter_last[29] ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[6] <= (((((((((((ethmac_crc32_inserter_last[30] ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]);
	ethmac_crc32_inserter_next[7] <= (((((((((ethmac_crc32_inserter_last[31] ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[8] <= ((((((((ethmac_crc32_inserter_last[0] ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_data1[6]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[9] <= ((((((((ethmac_crc32_inserter_last[1] ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_data1[6]);
	ethmac_crc32_inserter_next[10] <= ((((((((ethmac_crc32_inserter_last[2] ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[11] <= ((((((((ethmac_crc32_inserter_last[3] ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_data1[6]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[12] <= ((((((((((((ethmac_crc32_inserter_last[4] ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_data1[6]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[13] <= ((((((((((((ethmac_crc32_inserter_last[5] ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]);
	ethmac_crc32_inserter_next[14] <= ((((((((((ethmac_crc32_inserter_last[6] ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]);
	ethmac_crc32_inserter_next[15] <= ((((((((ethmac_crc32_inserter_last[7] ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]);
	ethmac_crc32_inserter_next[16] <= ((((((ethmac_crc32_inserter_last[8] ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[17] <= ((((((ethmac_crc32_inserter_last[9] ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_data1[6]);
	ethmac_crc32_inserter_next[18] <= ((((((ethmac_crc32_inserter_last[10] ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]);
	ethmac_crc32_inserter_next[19] <= ((((ethmac_crc32_inserter_last[11] ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]);
	ethmac_crc32_inserter_next[20] <= ((ethmac_crc32_inserter_last[12] ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]);
	ethmac_crc32_inserter_next[21] <= ((ethmac_crc32_inserter_last[13] ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]);
	ethmac_crc32_inserter_next[22] <= ((ethmac_crc32_inserter_last[14] ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[23] <= ((((((ethmac_crc32_inserter_last[15] ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_data1[6]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[24] <= ((((((ethmac_crc32_inserter_last[16] ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]);
	ethmac_crc32_inserter_next[25] <= ((((ethmac_crc32_inserter_last[17] ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]);
	ethmac_crc32_inserter_next[26] <= ((((((((ethmac_crc32_inserter_last[18] ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]) ^ ethmac_crc32_inserter_last[24]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_data1[7]);
	ethmac_crc32_inserter_next[27] <= ((((((((ethmac_crc32_inserter_last[19] ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]) ^ ethmac_crc32_inserter_last[25]) ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_data1[6]);
	ethmac_crc32_inserter_next[28] <= ((((((ethmac_crc32_inserter_last[20] ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]) ^ ethmac_crc32_inserter_last[26]) ^ ethmac_crc32_inserter_data1[5]);
	ethmac_crc32_inserter_next[29] <= ((((((ethmac_crc32_inserter_last[21] ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_last[30]) ^ ethmac_crc32_inserter_data1[1]) ^ ethmac_crc32_inserter_last[27]) ^ ethmac_crc32_inserter_data1[4]);
	ethmac_crc32_inserter_next[30] <= ((((ethmac_crc32_inserter_last[22] ^ ethmac_crc32_inserter_last[31]) ^ ethmac_crc32_inserter_data1[0]) ^ ethmac_crc32_inserter_last[28]) ^ ethmac_crc32_inserter_data1[3]);
	ethmac_crc32_inserter_next[31] <= ((ethmac_crc32_inserter_last[23] ^ ethmac_crc32_inserter_last[29]) ^ ethmac_crc32_inserter_data1[2]);
end
always @(*) begin
	ethmac_crc32_inserter_is_ongoing0 <= 1'd0;
	ethmac_crc32_inserter_sink_ready <= 1'd0;
	ethmac_crc32_inserter_is_ongoing1 <= 1'd0;
	ethmac_crc32_inserter_ce <= 1'd0;
	ethmac_crc32_inserter_reset <= 1'd0;
	ethmac_crc32_inserter_source_valid <= 1'd0;
	ethmac_crc32_inserter_source_first <= 1'd0;
	liteethmaccrc32inserter_next_state <= 2'd0;
	ethmac_crc32_inserter_source_last <= 1'd0;
	ethmac_crc32_inserter_source_payload_data <= 8'd0;
	ethmac_crc32_inserter_source_payload_last_be <= 1'd0;
	ethmac_crc32_inserter_source_payload_error <= 1'd0;
	ethmac_crc32_inserter_data0 <= 8'd0;
	liteethmaccrc32inserter_next_state <= liteethmaccrc32inserter_state;
	case (liteethmaccrc32inserter_state)
		1'd1: begin
			ethmac_crc32_inserter_ce <= (ethmac_crc32_inserter_sink_valid & ethmac_crc32_inserter_source_ready);
			ethmac_crc32_inserter_data0 <= ethmac_crc32_inserter_sink_payload_data;
			ethmac_crc32_inserter_source_valid <= ethmac_crc32_inserter_sink_valid;
			ethmac_crc32_inserter_sink_ready <= ethmac_crc32_inserter_source_ready;
			ethmac_crc32_inserter_source_first <= ethmac_crc32_inserter_sink_first;
			ethmac_crc32_inserter_source_last <= ethmac_crc32_inserter_sink_last;
			ethmac_crc32_inserter_source_payload_data <= ethmac_crc32_inserter_sink_payload_data;
			ethmac_crc32_inserter_source_payload_last_be <= ethmac_crc32_inserter_sink_payload_last_be;
			ethmac_crc32_inserter_source_payload_error <= ethmac_crc32_inserter_sink_payload_error;
			ethmac_crc32_inserter_source_last <= 1'd0;
			if (((ethmac_crc32_inserter_sink_valid & ethmac_crc32_inserter_sink_last) & ethmac_crc32_inserter_source_ready)) begin
				liteethmaccrc32inserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			ethmac_crc32_inserter_source_valid <= 1'd1;
			case (ethmac_crc32_inserter_cnt)
				1'd0: begin
					ethmac_crc32_inserter_source_payload_data <= ethmac_crc32_inserter_value[31:24];
				end
				1'd1: begin
					ethmac_crc32_inserter_source_payload_data <= ethmac_crc32_inserter_value[23:16];
				end
				2'd2: begin
					ethmac_crc32_inserter_source_payload_data <= ethmac_crc32_inserter_value[15:8];
				end
				default: begin
					ethmac_crc32_inserter_source_payload_data <= ethmac_crc32_inserter_value[7:0];
				end
			endcase
			if (ethmac_crc32_inserter_cnt_done) begin
				ethmac_crc32_inserter_source_last <= 1'd1;
				if (ethmac_crc32_inserter_source_ready) begin
					liteethmaccrc32inserter_next_state <= 1'd0;
				end
			end
			ethmac_crc32_inserter_is_ongoing1 <= 1'd1;
		end
		default: begin
			ethmac_crc32_inserter_reset <= 1'd1;
			ethmac_crc32_inserter_sink_ready <= 1'd1;
			if (ethmac_crc32_inserter_sink_valid) begin
				ethmac_crc32_inserter_sink_ready <= 1'd0;
				liteethmaccrc32inserter_next_state <= 1'd1;
			end
			ethmac_crc32_inserter_is_ongoing0 <= 1'd1;
		end
	endcase
end
assign ethmac_crc32_checker_fifo_full = (ethmac_crc32_checker_syncfifo_level == 3'd4);
assign ethmac_crc32_checker_fifo_in = (ethmac_crc32_checker_sink_sink_valid & ((~ethmac_crc32_checker_fifo_full) | ethmac_crc32_checker_fifo_out));
assign ethmac_crc32_checker_fifo_out = (ethmac_crc32_checker_source_source_valid & ethmac_crc32_checker_source_source_ready);
assign ethmac_crc32_checker_syncfifo_sink_first = ethmac_crc32_checker_sink_sink_first;
assign ethmac_crc32_checker_syncfifo_sink_last = ethmac_crc32_checker_sink_sink_last;
assign ethmac_crc32_checker_syncfifo_sink_payload_data = ethmac_crc32_checker_sink_sink_payload_data;
assign ethmac_crc32_checker_syncfifo_sink_payload_last_be = ethmac_crc32_checker_sink_sink_payload_last_be;
assign ethmac_crc32_checker_syncfifo_sink_payload_error = ethmac_crc32_checker_sink_sink_payload_error;
always @(*) begin
	ethmac_crc32_checker_syncfifo_sink_valid <= 1'd0;
	ethmac_crc32_checker_syncfifo_sink_valid <= ethmac_crc32_checker_sink_sink_valid;
	ethmac_crc32_checker_syncfifo_sink_valid <= ethmac_crc32_checker_fifo_in;
end
always @(*) begin
	ethmac_crc32_checker_sink_sink_ready <= 1'd0;
	ethmac_crc32_checker_sink_sink_ready <= ethmac_crc32_checker_syncfifo_sink_ready;
	ethmac_crc32_checker_sink_sink_ready <= ethmac_crc32_checker_fifo_in;
end
assign ethmac_crc32_checker_source_source_valid = (ethmac_crc32_checker_sink_sink_valid & ethmac_crc32_checker_fifo_full);
assign ethmac_crc32_checker_source_source_last = ethmac_crc32_checker_sink_sink_last;
assign ethmac_crc32_checker_syncfifo_source_ready = ethmac_crc32_checker_fifo_out;
assign ethmac_crc32_checker_source_source_payload_data = ethmac_crc32_checker_syncfifo_source_payload_data;
assign ethmac_crc32_checker_source_source_payload_last_be = ethmac_crc32_checker_syncfifo_source_payload_last_be;
always @(*) begin
	ethmac_crc32_checker_source_source_payload_error <= 1'd0;
	ethmac_crc32_checker_source_source_payload_error <= ethmac_crc32_checker_syncfifo_source_payload_error;
	ethmac_crc32_checker_source_source_payload_error <= (ethmac_crc32_checker_sink_sink_payload_error | ethmac_crc32_checker_crc_error);
end
assign ethmac_crc32_checker_error = ((ethmac_crc32_checker_source_source_valid & ethmac_crc32_checker_source_source_last) & ethmac_crc32_checker_crc_error);
assign ethmac_crc32_checker_crc_data0 = ethmac_crc32_checker_sink_sink_payload_data;
assign ethmac_crc32_checker_crc_data1 = ethmac_crc32_checker_crc_data0;
assign ethmac_crc32_checker_crc_last = ethmac_crc32_checker_crc_reg;
assign ethmac_crc32_checker_crc_value = (~{ethmac_crc32_checker_crc_reg[0], ethmac_crc32_checker_crc_reg[1], ethmac_crc32_checker_crc_reg[2], ethmac_crc32_checker_crc_reg[3], ethmac_crc32_checker_crc_reg[4], ethmac_crc32_checker_crc_reg[5], ethmac_crc32_checker_crc_reg[6], ethmac_crc32_checker_crc_reg[7], ethmac_crc32_checker_crc_reg[8], ethmac_crc32_checker_crc_reg[9], ethmac_crc32_checker_crc_reg[10], ethmac_crc32_checker_crc_reg[11], ethmac_crc32_checker_crc_reg[12], ethmac_crc32_checker_crc_reg[13], ethmac_crc32_checker_crc_reg[14], ethmac_crc32_checker_crc_reg[15], ethmac_crc32_checker_crc_reg[16], ethmac_crc32_checker_crc_reg[17], ethmac_crc32_checker_crc_reg[18], ethmac_crc32_checker_crc_reg[19], ethmac_crc32_checker_crc_reg[20], ethmac_crc32_checker_crc_reg[21], ethmac_crc32_checker_crc_reg[22], ethmac_crc32_checker_crc_reg[23], ethmac_crc32_checker_crc_reg[24], ethmac_crc32_checker_crc_reg[25], ethmac_crc32_checker_crc_reg[26], ethmac_crc32_checker_crc_reg[27], ethmac_crc32_checker_crc_reg[28], ethmac_crc32_checker_crc_reg[29], ethmac_crc32_checker_crc_reg[30], ethmac_crc32_checker_crc_reg[31]});
assign ethmac_crc32_checker_crc_error = (ethmac_crc32_checker_crc_next != 32'd3338984827);
always @(*) begin
	ethmac_crc32_checker_crc_next <= 32'd0;
	ethmac_crc32_checker_crc_next[0] <= (((ethmac_crc32_checker_crc_last[24] ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[1] <= (((((((ethmac_crc32_checker_crc_last[25] ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[2] <= (((((((((ethmac_crc32_checker_crc_last[26] ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[3] <= (((((((ethmac_crc32_checker_crc_last[27] ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]);
	ethmac_crc32_checker_crc_next[4] <= (((((((((ethmac_crc32_checker_crc_last[28] ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[5] <= (((((((((((((ethmac_crc32_checker_crc_last[29] ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[6] <= (((((((((((ethmac_crc32_checker_crc_last[30] ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]);
	ethmac_crc32_checker_crc_next[7] <= (((((((((ethmac_crc32_checker_crc_last[31] ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[8] <= ((((((((ethmac_crc32_checker_crc_last[0] ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_data1[6]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[9] <= ((((((((ethmac_crc32_checker_crc_last[1] ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_data1[6]);
	ethmac_crc32_checker_crc_next[10] <= ((((((((ethmac_crc32_checker_crc_last[2] ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[11] <= ((((((((ethmac_crc32_checker_crc_last[3] ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_data1[6]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[12] <= ((((((((((((ethmac_crc32_checker_crc_last[4] ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_data1[6]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[13] <= ((((((((((((ethmac_crc32_checker_crc_last[5] ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]);
	ethmac_crc32_checker_crc_next[14] <= ((((((((((ethmac_crc32_checker_crc_last[6] ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]);
	ethmac_crc32_checker_crc_next[15] <= ((((((((ethmac_crc32_checker_crc_last[7] ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]);
	ethmac_crc32_checker_crc_next[16] <= ((((((ethmac_crc32_checker_crc_last[8] ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[17] <= ((((((ethmac_crc32_checker_crc_last[9] ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_data1[6]);
	ethmac_crc32_checker_crc_next[18] <= ((((((ethmac_crc32_checker_crc_last[10] ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]);
	ethmac_crc32_checker_crc_next[19] <= ((((ethmac_crc32_checker_crc_last[11] ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]);
	ethmac_crc32_checker_crc_next[20] <= ((ethmac_crc32_checker_crc_last[12] ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]);
	ethmac_crc32_checker_crc_next[21] <= ((ethmac_crc32_checker_crc_last[13] ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]);
	ethmac_crc32_checker_crc_next[22] <= ((ethmac_crc32_checker_crc_last[14] ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[23] <= ((((((ethmac_crc32_checker_crc_last[15] ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_data1[6]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[24] <= ((((((ethmac_crc32_checker_crc_last[16] ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]);
	ethmac_crc32_checker_crc_next[25] <= ((((ethmac_crc32_checker_crc_last[17] ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]);
	ethmac_crc32_checker_crc_next[26] <= ((((((((ethmac_crc32_checker_crc_last[18] ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]) ^ ethmac_crc32_checker_crc_last[24]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_data1[7]);
	ethmac_crc32_checker_crc_next[27] <= ((((((((ethmac_crc32_checker_crc_last[19] ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]) ^ ethmac_crc32_checker_crc_last[25]) ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_data1[6]);
	ethmac_crc32_checker_crc_next[28] <= ((((((ethmac_crc32_checker_crc_last[20] ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]) ^ ethmac_crc32_checker_crc_last[26]) ^ ethmac_crc32_checker_crc_data1[5]);
	ethmac_crc32_checker_crc_next[29] <= ((((((ethmac_crc32_checker_crc_last[21] ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_last[30]) ^ ethmac_crc32_checker_crc_data1[1]) ^ ethmac_crc32_checker_crc_last[27]) ^ ethmac_crc32_checker_crc_data1[4]);
	ethmac_crc32_checker_crc_next[30] <= ((((ethmac_crc32_checker_crc_last[22] ^ ethmac_crc32_checker_crc_last[31]) ^ ethmac_crc32_checker_crc_data1[0]) ^ ethmac_crc32_checker_crc_last[28]) ^ ethmac_crc32_checker_crc_data1[3]);
	ethmac_crc32_checker_crc_next[31] <= ((ethmac_crc32_checker_crc_last[23] ^ ethmac_crc32_checker_crc_last[29]) ^ ethmac_crc32_checker_crc_data1[2]);
end
assign ethmac_crc32_checker_syncfifo_syncfifo_din = {ethmac_crc32_checker_syncfifo_fifo_in_last, ethmac_crc32_checker_syncfifo_fifo_in_first, ethmac_crc32_checker_syncfifo_fifo_in_payload_error, ethmac_crc32_checker_syncfifo_fifo_in_payload_last_be, ethmac_crc32_checker_syncfifo_fifo_in_payload_data};
assign {ethmac_crc32_checker_syncfifo_fifo_out_last, ethmac_crc32_checker_syncfifo_fifo_out_first, ethmac_crc32_checker_syncfifo_fifo_out_payload_error, ethmac_crc32_checker_syncfifo_fifo_out_payload_last_be, ethmac_crc32_checker_syncfifo_fifo_out_payload_data} = ethmac_crc32_checker_syncfifo_syncfifo_dout;
assign ethmac_crc32_checker_syncfifo_sink_ready = ethmac_crc32_checker_syncfifo_syncfifo_writable;
assign ethmac_crc32_checker_syncfifo_syncfifo_we = ethmac_crc32_checker_syncfifo_sink_valid;
assign ethmac_crc32_checker_syncfifo_fifo_in_first = ethmac_crc32_checker_syncfifo_sink_first;
assign ethmac_crc32_checker_syncfifo_fifo_in_last = ethmac_crc32_checker_syncfifo_sink_last;
assign ethmac_crc32_checker_syncfifo_fifo_in_payload_data = ethmac_crc32_checker_syncfifo_sink_payload_data;
assign ethmac_crc32_checker_syncfifo_fifo_in_payload_last_be = ethmac_crc32_checker_syncfifo_sink_payload_last_be;
assign ethmac_crc32_checker_syncfifo_fifo_in_payload_error = ethmac_crc32_checker_syncfifo_sink_payload_error;
assign ethmac_crc32_checker_syncfifo_source_valid = ethmac_crc32_checker_syncfifo_syncfifo_readable;
assign ethmac_crc32_checker_syncfifo_source_first = ethmac_crc32_checker_syncfifo_fifo_out_first;
assign ethmac_crc32_checker_syncfifo_source_last = ethmac_crc32_checker_syncfifo_fifo_out_last;
assign ethmac_crc32_checker_syncfifo_source_payload_data = ethmac_crc32_checker_syncfifo_fifo_out_payload_data;
assign ethmac_crc32_checker_syncfifo_source_payload_last_be = ethmac_crc32_checker_syncfifo_fifo_out_payload_last_be;
assign ethmac_crc32_checker_syncfifo_source_payload_error = ethmac_crc32_checker_syncfifo_fifo_out_payload_error;
assign ethmac_crc32_checker_syncfifo_syncfifo_re = ethmac_crc32_checker_syncfifo_source_ready;
always @(*) begin
	ethmac_crc32_checker_syncfifo_wrport_adr <= 3'd0;
	if (ethmac_crc32_checker_syncfifo_replace) begin
		ethmac_crc32_checker_syncfifo_wrport_adr <= (ethmac_crc32_checker_syncfifo_produce - 1'd1);
	end else begin
		ethmac_crc32_checker_syncfifo_wrport_adr <= ethmac_crc32_checker_syncfifo_produce;
	end
end
assign ethmac_crc32_checker_syncfifo_wrport_dat_w = ethmac_crc32_checker_syncfifo_syncfifo_din;
assign ethmac_crc32_checker_syncfifo_wrport_we = (ethmac_crc32_checker_syncfifo_syncfifo_we & (ethmac_crc32_checker_syncfifo_syncfifo_writable | ethmac_crc32_checker_syncfifo_replace));
assign ethmac_crc32_checker_syncfifo_do_read = (ethmac_crc32_checker_syncfifo_syncfifo_readable & ethmac_crc32_checker_syncfifo_syncfifo_re);
assign ethmac_crc32_checker_syncfifo_rdport_adr = ethmac_crc32_checker_syncfifo_consume;
assign ethmac_crc32_checker_syncfifo_syncfifo_dout = ethmac_crc32_checker_syncfifo_rdport_dat_r;
assign ethmac_crc32_checker_syncfifo_syncfifo_writable = (ethmac_crc32_checker_syncfifo_level != 3'd5);
assign ethmac_crc32_checker_syncfifo_syncfifo_readable = (ethmac_crc32_checker_syncfifo_level != 1'd0);
always @(*) begin
	liteethmaccrc32checker_next_state <= 2'd0;
	ethmac_crc32_checker_crc_ce <= 1'd0;
	ethmac_crc32_checker_crc_reset <= 1'd0;
	ethmac_crc32_checker_fifo_reset <= 1'd0;
	liteethmaccrc32checker_next_state <= liteethmaccrc32checker_state;
	case (liteethmaccrc32checker_state)
		1'd1: begin
			if ((ethmac_crc32_checker_sink_sink_valid & ethmac_crc32_checker_sink_sink_ready)) begin
				ethmac_crc32_checker_crc_ce <= 1'd1;
				liteethmaccrc32checker_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((ethmac_crc32_checker_sink_sink_valid & ethmac_crc32_checker_sink_sink_ready)) begin
				ethmac_crc32_checker_crc_ce <= 1'd1;
				if (ethmac_crc32_checker_sink_sink_last) begin
					liteethmaccrc32checker_next_state <= 1'd0;
				end
			end
		end
		default: begin
			ethmac_crc32_checker_crc_reset <= 1'd1;
			ethmac_crc32_checker_fifo_reset <= 1'd1;
			liteethmaccrc32checker_next_state <= 1'd1;
		end
	endcase
end
assign ethmac_ps_preamble_error_o = (ethmac_ps_preamble_error_toggle_o ^ ethmac_ps_preamble_error_toggle_o_r);
assign ethmac_ps_crc_error_o = (ethmac_ps_crc_error_toggle_o ^ ethmac_ps_crc_error_toggle_o_r);
assign ethmac_padding_inserter_counter_done = (ethmac_padding_inserter_counter >= 6'd59);
always @(*) begin
	ethmac_padding_inserter_counter_reset <= 1'd0;
	ethmac_padding_inserter_counter_ce <= 1'd0;
	ethmac_padding_inserter_sink_ready <= 1'd0;
	ethmac_padding_inserter_source_valid <= 1'd0;
	ethmac_padding_inserter_source_first <= 1'd0;
	liteethmacpaddinginserter_next_state <= 1'd0;
	ethmac_padding_inserter_source_last <= 1'd0;
	ethmac_padding_inserter_source_payload_data <= 8'd0;
	ethmac_padding_inserter_source_payload_last_be <= 1'd0;
	ethmac_padding_inserter_source_payload_error <= 1'd0;
	liteethmacpaddinginserter_next_state <= liteethmacpaddinginserter_state;
	case (liteethmacpaddinginserter_state)
		1'd1: begin
			ethmac_padding_inserter_source_valid <= 1'd1;
			ethmac_padding_inserter_source_last <= ethmac_padding_inserter_counter_done;
			ethmac_padding_inserter_source_payload_data <= 1'd0;
			if ((ethmac_padding_inserter_source_valid & ethmac_padding_inserter_source_ready)) begin
				ethmac_padding_inserter_counter_ce <= 1'd1;
				if (ethmac_padding_inserter_counter_done) begin
					ethmac_padding_inserter_counter_reset <= 1'd1;
					liteethmacpaddinginserter_next_state <= 1'd0;
				end
			end
		end
		default: begin
			ethmac_padding_inserter_source_valid <= ethmac_padding_inserter_sink_valid;
			ethmac_padding_inserter_sink_ready <= ethmac_padding_inserter_source_ready;
			ethmac_padding_inserter_source_first <= ethmac_padding_inserter_sink_first;
			ethmac_padding_inserter_source_last <= ethmac_padding_inserter_sink_last;
			ethmac_padding_inserter_source_payload_data <= ethmac_padding_inserter_sink_payload_data;
			ethmac_padding_inserter_source_payload_last_be <= ethmac_padding_inserter_sink_payload_last_be;
			ethmac_padding_inserter_source_payload_error <= ethmac_padding_inserter_sink_payload_error;
			if ((ethmac_padding_inserter_source_valid & ethmac_padding_inserter_source_ready)) begin
				ethmac_padding_inserter_counter_ce <= 1'd1;
				if (ethmac_padding_inserter_sink_last) begin
					if ((~ethmac_padding_inserter_counter_done)) begin
						ethmac_padding_inserter_source_last <= 1'd0;
						liteethmacpaddinginserter_next_state <= 1'd1;
					end else begin
						ethmac_padding_inserter_counter_reset <= 1'd1;
					end
				end
			end
		end
	endcase
end
assign ethmac_padding_checker_source_valid = ethmac_padding_checker_sink_valid;
assign ethmac_padding_checker_sink_ready = ethmac_padding_checker_source_ready;
assign ethmac_padding_checker_source_first = ethmac_padding_checker_sink_first;
assign ethmac_padding_checker_source_last = ethmac_padding_checker_sink_last;
assign ethmac_padding_checker_source_payload_data = ethmac_padding_checker_sink_payload_data;
assign ethmac_padding_checker_source_payload_last_be = ethmac_padding_checker_sink_payload_last_be;
assign ethmac_padding_checker_source_payload_error = ethmac_padding_checker_sink_payload_error;
assign ethmac_tx_last_be_source_valid = (ethmac_tx_last_be_sink_valid & ethmac_tx_last_be_ongoing);
assign ethmac_tx_last_be_source_last = ethmac_tx_last_be_sink_payload_last_be;
assign ethmac_tx_last_be_source_payload_data = ethmac_tx_last_be_sink_payload_data;
assign ethmac_tx_last_be_sink_ready = ethmac_tx_last_be_source_ready;
assign ethmac_rx_last_be_source_valid = ethmac_rx_last_be_sink_valid;
assign ethmac_rx_last_be_sink_ready = ethmac_rx_last_be_source_ready;
assign ethmac_rx_last_be_source_first = ethmac_rx_last_be_sink_first;
assign ethmac_rx_last_be_source_last = ethmac_rx_last_be_sink_last;
assign ethmac_rx_last_be_source_payload_data = ethmac_rx_last_be_sink_payload_data;
assign ethmac_rx_last_be_source_payload_error = ethmac_rx_last_be_sink_payload_error;
always @(*) begin
	ethmac_rx_last_be_source_payload_last_be <= 1'd0;
	ethmac_rx_last_be_source_payload_last_be <= ethmac_rx_last_be_sink_payload_last_be;
	ethmac_rx_last_be_source_payload_last_be <= ethmac_rx_last_be_sink_last;
end
assign ethmac_tx_converter_converter_sink_valid = ethmac_tx_converter_sink_valid;
assign ethmac_tx_converter_converter_sink_first = ethmac_tx_converter_sink_first;
assign ethmac_tx_converter_converter_sink_last = ethmac_tx_converter_sink_last;
assign ethmac_tx_converter_sink_ready = ethmac_tx_converter_converter_sink_ready;
always @(*) begin
	ethmac_tx_converter_converter_sink_payload_data <= 40'd0;
	ethmac_tx_converter_converter_sink_payload_data[7:0] <= ethmac_tx_converter_sink_payload_data[7:0];
	ethmac_tx_converter_converter_sink_payload_data[8] <= ethmac_tx_converter_sink_payload_last_be[0];
	ethmac_tx_converter_converter_sink_payload_data[9] <= ethmac_tx_converter_sink_payload_error[0];
	ethmac_tx_converter_converter_sink_payload_data[17:10] <= ethmac_tx_converter_sink_payload_data[15:8];
	ethmac_tx_converter_converter_sink_payload_data[18] <= ethmac_tx_converter_sink_payload_last_be[1];
	ethmac_tx_converter_converter_sink_payload_data[19] <= ethmac_tx_converter_sink_payload_error[1];
	ethmac_tx_converter_converter_sink_payload_data[27:20] <= ethmac_tx_converter_sink_payload_data[23:16];
	ethmac_tx_converter_converter_sink_payload_data[28] <= ethmac_tx_converter_sink_payload_last_be[2];
	ethmac_tx_converter_converter_sink_payload_data[29] <= ethmac_tx_converter_sink_payload_error[2];
	ethmac_tx_converter_converter_sink_payload_data[37:30] <= ethmac_tx_converter_sink_payload_data[31:24];
	ethmac_tx_converter_converter_sink_payload_data[38] <= ethmac_tx_converter_sink_payload_last_be[3];
	ethmac_tx_converter_converter_sink_payload_data[39] <= ethmac_tx_converter_sink_payload_error[3];
end
assign ethmac_tx_converter_source_valid = ethmac_tx_converter_source_source_valid;
assign ethmac_tx_converter_source_first = ethmac_tx_converter_source_source_first;
assign ethmac_tx_converter_source_last = ethmac_tx_converter_source_source_last;
assign ethmac_tx_converter_source_source_ready = ethmac_tx_converter_source_ready;
assign {ethmac_tx_converter_source_payload_error, ethmac_tx_converter_source_payload_last_be, ethmac_tx_converter_source_payload_data} = ethmac_tx_converter_source_source_payload_data;
assign ethmac_tx_converter_source_source_valid = ethmac_tx_converter_converter_source_valid;
assign ethmac_tx_converter_converter_source_ready = ethmac_tx_converter_source_source_ready;
assign ethmac_tx_converter_source_source_first = ethmac_tx_converter_converter_source_first;
assign ethmac_tx_converter_source_source_last = ethmac_tx_converter_converter_source_last;
assign ethmac_tx_converter_source_source_payload_data = ethmac_tx_converter_converter_source_payload_data;
assign ethmac_tx_converter_converter_first = (ethmac_tx_converter_converter_mux == 1'd0);
assign ethmac_tx_converter_converter_last = (ethmac_tx_converter_converter_mux == 2'd3);
assign ethmac_tx_converter_converter_source_valid = ethmac_tx_converter_converter_sink_valid;
assign ethmac_tx_converter_converter_source_first = (ethmac_tx_converter_converter_sink_first & ethmac_tx_converter_converter_first);
assign ethmac_tx_converter_converter_source_last = (ethmac_tx_converter_converter_sink_last & ethmac_tx_converter_converter_last);
assign ethmac_tx_converter_converter_sink_ready = (ethmac_tx_converter_converter_last & ethmac_tx_converter_converter_source_ready);
always @(*) begin
	ethmac_tx_converter_converter_source_payload_data <= 10'd0;
	case (ethmac_tx_converter_converter_mux)
		1'd0: begin
			ethmac_tx_converter_converter_source_payload_data <= ethmac_tx_converter_converter_sink_payload_data[39:30];
		end
		1'd1: begin
			ethmac_tx_converter_converter_source_payload_data <= ethmac_tx_converter_converter_sink_payload_data[29:20];
		end
		2'd2: begin
			ethmac_tx_converter_converter_source_payload_data <= ethmac_tx_converter_converter_sink_payload_data[19:10];
		end
		default: begin
			ethmac_tx_converter_converter_source_payload_data <= ethmac_tx_converter_converter_sink_payload_data[9:0];
		end
	endcase
end
assign ethmac_tx_converter_converter_source_payload_valid_token_count = ethmac_tx_converter_converter_last;
assign ethmac_rx_converter_converter_sink_valid = ethmac_rx_converter_sink_valid;
assign ethmac_rx_converter_converter_sink_first = ethmac_rx_converter_sink_first;
assign ethmac_rx_converter_converter_sink_last = ethmac_rx_converter_sink_last;
assign ethmac_rx_converter_sink_ready = ethmac_rx_converter_converter_sink_ready;
assign ethmac_rx_converter_converter_sink_payload_data = {ethmac_rx_converter_sink_payload_error, ethmac_rx_converter_sink_payload_last_be, ethmac_rx_converter_sink_payload_data};
assign ethmac_rx_converter_source_valid = ethmac_rx_converter_source_source_valid;
assign ethmac_rx_converter_source_first = ethmac_rx_converter_source_source_first;
assign ethmac_rx_converter_source_last = ethmac_rx_converter_source_source_last;
assign ethmac_rx_converter_source_source_ready = ethmac_rx_converter_source_ready;
always @(*) begin
	ethmac_rx_converter_source_payload_data <= 32'd0;
	ethmac_rx_converter_source_payload_data[7:0] <= ethmac_rx_converter_source_source_payload_data[7:0];
	ethmac_rx_converter_source_payload_data[15:8] <= ethmac_rx_converter_source_source_payload_data[17:10];
	ethmac_rx_converter_source_payload_data[23:16] <= ethmac_rx_converter_source_source_payload_data[27:20];
	ethmac_rx_converter_source_payload_data[31:24] <= ethmac_rx_converter_source_source_payload_data[37:30];
end
always @(*) begin
	ethmac_rx_converter_source_payload_last_be <= 4'd0;
	ethmac_rx_converter_source_payload_last_be[0] <= ethmac_rx_converter_source_source_payload_data[8];
	ethmac_rx_converter_source_payload_last_be[1] <= ethmac_rx_converter_source_source_payload_data[18];
	ethmac_rx_converter_source_payload_last_be[2] <= ethmac_rx_converter_source_source_payload_data[28];
	ethmac_rx_converter_source_payload_last_be[3] <= ethmac_rx_converter_source_source_payload_data[38];
end
always @(*) begin
	ethmac_rx_converter_source_payload_error <= 4'd0;
	ethmac_rx_converter_source_payload_error[0] <= ethmac_rx_converter_source_source_payload_data[9];
	ethmac_rx_converter_source_payload_error[1] <= ethmac_rx_converter_source_source_payload_data[19];
	ethmac_rx_converter_source_payload_error[2] <= ethmac_rx_converter_source_source_payload_data[29];
	ethmac_rx_converter_source_payload_error[3] <= ethmac_rx_converter_source_source_payload_data[39];
end
assign ethmac_rx_converter_source_source_valid = ethmac_rx_converter_converter_source_valid;
assign ethmac_rx_converter_converter_source_ready = ethmac_rx_converter_source_source_ready;
assign ethmac_rx_converter_source_source_first = ethmac_rx_converter_converter_source_first;
assign ethmac_rx_converter_source_source_last = ethmac_rx_converter_converter_source_last;
assign ethmac_rx_converter_source_source_payload_data = ethmac_rx_converter_converter_source_payload_data;
assign ethmac_rx_converter_converter_sink_ready = ((~ethmac_rx_converter_converter_strobe_all) | ethmac_rx_converter_converter_source_ready);
assign ethmac_rx_converter_converter_source_valid = ethmac_rx_converter_converter_strobe_all;
assign ethmac_rx_converter_converter_load_part = (ethmac_rx_converter_converter_sink_valid & ethmac_rx_converter_converter_sink_ready);
assign ethmac_tx_cdc_asyncfifo_din = {ethmac_tx_cdc_fifo_in_last, ethmac_tx_cdc_fifo_in_first, ethmac_tx_cdc_fifo_in_payload_error, ethmac_tx_cdc_fifo_in_payload_last_be, ethmac_tx_cdc_fifo_in_payload_data};
assign {ethmac_tx_cdc_fifo_out_last, ethmac_tx_cdc_fifo_out_first, ethmac_tx_cdc_fifo_out_payload_error, ethmac_tx_cdc_fifo_out_payload_last_be, ethmac_tx_cdc_fifo_out_payload_data} = ethmac_tx_cdc_asyncfifo_dout;
assign ethmac_tx_cdc_sink_ready = ethmac_tx_cdc_asyncfifo_writable;
assign ethmac_tx_cdc_asyncfifo_we = ethmac_tx_cdc_sink_valid;
assign ethmac_tx_cdc_fifo_in_first = ethmac_tx_cdc_sink_first;
assign ethmac_tx_cdc_fifo_in_last = ethmac_tx_cdc_sink_last;
assign ethmac_tx_cdc_fifo_in_payload_data = ethmac_tx_cdc_sink_payload_data;
assign ethmac_tx_cdc_fifo_in_payload_last_be = ethmac_tx_cdc_sink_payload_last_be;
assign ethmac_tx_cdc_fifo_in_payload_error = ethmac_tx_cdc_sink_payload_error;
assign ethmac_tx_cdc_source_valid = ethmac_tx_cdc_asyncfifo_readable;
assign ethmac_tx_cdc_source_first = ethmac_tx_cdc_fifo_out_first;
assign ethmac_tx_cdc_source_last = ethmac_tx_cdc_fifo_out_last;
assign ethmac_tx_cdc_source_payload_data = ethmac_tx_cdc_fifo_out_payload_data;
assign ethmac_tx_cdc_source_payload_last_be = ethmac_tx_cdc_fifo_out_payload_last_be;
assign ethmac_tx_cdc_source_payload_error = ethmac_tx_cdc_fifo_out_payload_error;
assign ethmac_tx_cdc_asyncfifo_re = ethmac_tx_cdc_source_ready;
assign ethmac_tx_cdc_graycounter0_ce = (ethmac_tx_cdc_asyncfifo_writable & ethmac_tx_cdc_asyncfifo_we);
assign ethmac_tx_cdc_graycounter1_ce = (ethmac_tx_cdc_asyncfifo_readable & ethmac_tx_cdc_asyncfifo_re);
assign ethmac_tx_cdc_asyncfifo_writable = (((ethmac_tx_cdc_graycounter0_q[6] == ethmac_tx_cdc_consume_wdomain[6]) | (ethmac_tx_cdc_graycounter0_q[5] == ethmac_tx_cdc_consume_wdomain[5])) | (ethmac_tx_cdc_graycounter0_q[4:0] != ethmac_tx_cdc_consume_wdomain[4:0]));
assign ethmac_tx_cdc_asyncfifo_readable = (ethmac_tx_cdc_graycounter1_q != ethmac_tx_cdc_produce_rdomain);
assign ethmac_tx_cdc_wrport_adr = ethmac_tx_cdc_graycounter0_q_binary[5:0];
assign ethmac_tx_cdc_wrport_dat_w = ethmac_tx_cdc_asyncfifo_din;
assign ethmac_tx_cdc_wrport_we = ethmac_tx_cdc_graycounter0_ce;
assign ethmac_tx_cdc_rdport_adr = ethmac_tx_cdc_graycounter1_q_next_binary[5:0];
assign ethmac_tx_cdc_asyncfifo_dout = ethmac_tx_cdc_rdport_dat_r;
always @(*) begin
	ethmac_tx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (ethmac_tx_cdc_graycounter0_ce) begin
		ethmac_tx_cdc_graycounter0_q_next_binary <= (ethmac_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		ethmac_tx_cdc_graycounter0_q_next_binary <= ethmac_tx_cdc_graycounter0_q_binary;
	end
end
assign ethmac_tx_cdc_graycounter0_q_next = (ethmac_tx_cdc_graycounter0_q_next_binary ^ ethmac_tx_cdc_graycounter0_q_next_binary[6:1]);
always @(*) begin
	ethmac_tx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (ethmac_tx_cdc_graycounter1_ce) begin
		ethmac_tx_cdc_graycounter1_q_next_binary <= (ethmac_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		ethmac_tx_cdc_graycounter1_q_next_binary <= ethmac_tx_cdc_graycounter1_q_binary;
	end
end
assign ethmac_tx_cdc_graycounter1_q_next = (ethmac_tx_cdc_graycounter1_q_next_binary ^ ethmac_tx_cdc_graycounter1_q_next_binary[6:1]);
assign ethmac_rx_cdc_asyncfifo_din = {ethmac_rx_cdc_fifo_in_last, ethmac_rx_cdc_fifo_in_first, ethmac_rx_cdc_fifo_in_payload_error, ethmac_rx_cdc_fifo_in_payload_last_be, ethmac_rx_cdc_fifo_in_payload_data};
assign {ethmac_rx_cdc_fifo_out_last, ethmac_rx_cdc_fifo_out_first, ethmac_rx_cdc_fifo_out_payload_error, ethmac_rx_cdc_fifo_out_payload_last_be, ethmac_rx_cdc_fifo_out_payload_data} = ethmac_rx_cdc_asyncfifo_dout;
assign ethmac_rx_cdc_sink_ready = ethmac_rx_cdc_asyncfifo_writable;
assign ethmac_rx_cdc_asyncfifo_we = ethmac_rx_cdc_sink_valid;
assign ethmac_rx_cdc_fifo_in_first = ethmac_rx_cdc_sink_first;
assign ethmac_rx_cdc_fifo_in_last = ethmac_rx_cdc_sink_last;
assign ethmac_rx_cdc_fifo_in_payload_data = ethmac_rx_cdc_sink_payload_data;
assign ethmac_rx_cdc_fifo_in_payload_last_be = ethmac_rx_cdc_sink_payload_last_be;
assign ethmac_rx_cdc_fifo_in_payload_error = ethmac_rx_cdc_sink_payload_error;
assign ethmac_rx_cdc_source_valid = ethmac_rx_cdc_asyncfifo_readable;
assign ethmac_rx_cdc_source_first = ethmac_rx_cdc_fifo_out_first;
assign ethmac_rx_cdc_source_last = ethmac_rx_cdc_fifo_out_last;
assign ethmac_rx_cdc_source_payload_data = ethmac_rx_cdc_fifo_out_payload_data;
assign ethmac_rx_cdc_source_payload_last_be = ethmac_rx_cdc_fifo_out_payload_last_be;
assign ethmac_rx_cdc_source_payload_error = ethmac_rx_cdc_fifo_out_payload_error;
assign ethmac_rx_cdc_asyncfifo_re = ethmac_rx_cdc_source_ready;
assign ethmac_rx_cdc_graycounter0_ce = (ethmac_rx_cdc_asyncfifo_writable & ethmac_rx_cdc_asyncfifo_we);
assign ethmac_rx_cdc_graycounter1_ce = (ethmac_rx_cdc_asyncfifo_readable & ethmac_rx_cdc_asyncfifo_re);
assign ethmac_rx_cdc_asyncfifo_writable = (((ethmac_rx_cdc_graycounter0_q[6] == ethmac_rx_cdc_consume_wdomain[6]) | (ethmac_rx_cdc_graycounter0_q[5] == ethmac_rx_cdc_consume_wdomain[5])) | (ethmac_rx_cdc_graycounter0_q[4:0] != ethmac_rx_cdc_consume_wdomain[4:0]));
assign ethmac_rx_cdc_asyncfifo_readable = (ethmac_rx_cdc_graycounter1_q != ethmac_rx_cdc_produce_rdomain);
assign ethmac_rx_cdc_wrport_adr = ethmac_rx_cdc_graycounter0_q_binary[5:0];
assign ethmac_rx_cdc_wrport_dat_w = ethmac_rx_cdc_asyncfifo_din;
assign ethmac_rx_cdc_wrport_we = ethmac_rx_cdc_graycounter0_ce;
assign ethmac_rx_cdc_rdport_adr = ethmac_rx_cdc_graycounter1_q_next_binary[5:0];
assign ethmac_rx_cdc_asyncfifo_dout = ethmac_rx_cdc_rdport_dat_r;
always @(*) begin
	ethmac_rx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (ethmac_rx_cdc_graycounter0_ce) begin
		ethmac_rx_cdc_graycounter0_q_next_binary <= (ethmac_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		ethmac_rx_cdc_graycounter0_q_next_binary <= ethmac_rx_cdc_graycounter0_q_binary;
	end
end
assign ethmac_rx_cdc_graycounter0_q_next = (ethmac_rx_cdc_graycounter0_q_next_binary ^ ethmac_rx_cdc_graycounter0_q_next_binary[6:1]);
always @(*) begin
	ethmac_rx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (ethmac_rx_cdc_graycounter1_ce) begin
		ethmac_rx_cdc_graycounter1_q_next_binary <= (ethmac_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		ethmac_rx_cdc_graycounter1_q_next_binary <= ethmac_rx_cdc_graycounter1_q_binary;
	end
end
assign ethmac_rx_cdc_graycounter1_q_next = (ethmac_rx_cdc_graycounter1_q_next_binary ^ ethmac_rx_cdc_graycounter1_q_next_binary[6:1]);
assign ethmac_tx_converter_sink_valid = ethmac_tx_cdc_source_valid;
assign ethmac_tx_cdc_source_ready = ethmac_tx_converter_sink_ready;
assign ethmac_tx_converter_sink_first = ethmac_tx_cdc_source_first;
assign ethmac_tx_converter_sink_last = ethmac_tx_cdc_source_last;
assign ethmac_tx_converter_sink_payload_data = ethmac_tx_cdc_source_payload_data;
assign ethmac_tx_converter_sink_payload_last_be = ethmac_tx_cdc_source_payload_last_be;
assign ethmac_tx_converter_sink_payload_error = ethmac_tx_cdc_source_payload_error;
assign ethmac_tx_last_be_sink_valid = ethmac_tx_converter_source_valid;
assign ethmac_tx_converter_source_ready = ethmac_tx_last_be_sink_ready;
assign ethmac_tx_last_be_sink_first = ethmac_tx_converter_source_first;
assign ethmac_tx_last_be_sink_last = ethmac_tx_converter_source_last;
assign ethmac_tx_last_be_sink_payload_data = ethmac_tx_converter_source_payload_data;
assign ethmac_tx_last_be_sink_payload_last_be = ethmac_tx_converter_source_payload_last_be;
assign ethmac_tx_last_be_sink_payload_error = ethmac_tx_converter_source_payload_error;
assign ethmac_padding_inserter_sink_valid = ethmac_tx_last_be_source_valid;
assign ethmac_tx_last_be_source_ready = ethmac_padding_inserter_sink_ready;
assign ethmac_padding_inserter_sink_first = ethmac_tx_last_be_source_first;
assign ethmac_padding_inserter_sink_last = ethmac_tx_last_be_source_last;
assign ethmac_padding_inserter_sink_payload_data = ethmac_tx_last_be_source_payload_data;
assign ethmac_padding_inserter_sink_payload_last_be = ethmac_tx_last_be_source_payload_last_be;
assign ethmac_padding_inserter_sink_payload_error = ethmac_tx_last_be_source_payload_error;
assign ethmac_crc32_inserter_sink_valid = ethmac_padding_inserter_source_valid;
assign ethmac_padding_inserter_source_ready = ethmac_crc32_inserter_sink_ready;
assign ethmac_crc32_inserter_sink_first = ethmac_padding_inserter_source_first;
assign ethmac_crc32_inserter_sink_last = ethmac_padding_inserter_source_last;
assign ethmac_crc32_inserter_sink_payload_data = ethmac_padding_inserter_source_payload_data;
assign ethmac_crc32_inserter_sink_payload_last_be = ethmac_padding_inserter_source_payload_last_be;
assign ethmac_crc32_inserter_sink_payload_error = ethmac_padding_inserter_source_payload_error;
assign ethmac_preamble_inserter_sink_valid = ethmac_crc32_inserter_source_valid;
assign ethmac_crc32_inserter_source_ready = ethmac_preamble_inserter_sink_ready;
assign ethmac_preamble_inserter_sink_first = ethmac_crc32_inserter_source_first;
assign ethmac_preamble_inserter_sink_last = ethmac_crc32_inserter_source_last;
assign ethmac_preamble_inserter_sink_payload_data = ethmac_crc32_inserter_source_payload_data;
assign ethmac_preamble_inserter_sink_payload_last_be = ethmac_crc32_inserter_source_payload_last_be;
assign ethmac_preamble_inserter_sink_payload_error = ethmac_crc32_inserter_source_payload_error;
assign ethmac_tx_gap_inserter_sink_valid = ethmac_preamble_inserter_source_valid;
assign ethmac_preamble_inserter_source_ready = ethmac_tx_gap_inserter_sink_ready;
assign ethmac_tx_gap_inserter_sink_first = ethmac_preamble_inserter_source_first;
assign ethmac_tx_gap_inserter_sink_last = ethmac_preamble_inserter_source_last;
assign ethmac_tx_gap_inserter_sink_payload_data = ethmac_preamble_inserter_source_payload_data;
assign ethmac_tx_gap_inserter_sink_payload_last_be = ethmac_preamble_inserter_source_payload_last_be;
assign ethmac_tx_gap_inserter_sink_payload_error = ethmac_preamble_inserter_source_payload_error;
assign ethphy_sink_valid = ethmac_tx_gap_inserter_source_valid;
assign ethmac_tx_gap_inserter_source_ready = ethphy_sink_ready;
assign ethphy_sink_first = ethmac_tx_gap_inserter_source_first;
assign ethphy_sink_last = ethmac_tx_gap_inserter_source_last;
assign ethphy_sink_payload_data = ethmac_tx_gap_inserter_source_payload_data;
assign ethphy_sink_payload_last_be = ethmac_tx_gap_inserter_source_payload_last_be;
assign ethphy_sink_payload_error = ethmac_tx_gap_inserter_source_payload_error;
assign ethmac_preamble_checker_sink_valid = ethphy_source_valid;
assign ethphy_source_ready = ethmac_preamble_checker_sink_ready;
assign ethmac_preamble_checker_sink_first = ethphy_source_first;
assign ethmac_preamble_checker_sink_last = ethphy_source_last;
assign ethmac_preamble_checker_sink_payload_data = ethphy_source_payload_data;
assign ethmac_preamble_checker_sink_payload_last_be = ethphy_source_payload_last_be;
assign ethmac_preamble_checker_sink_payload_error = ethphy_source_payload_error;
assign ethmac_crc32_checker_sink_sink_valid = ethmac_preamble_checker_source_valid;
assign ethmac_preamble_checker_source_ready = ethmac_crc32_checker_sink_sink_ready;
assign ethmac_crc32_checker_sink_sink_first = ethmac_preamble_checker_source_first;
assign ethmac_crc32_checker_sink_sink_last = ethmac_preamble_checker_source_last;
assign ethmac_crc32_checker_sink_sink_payload_data = ethmac_preamble_checker_source_payload_data;
assign ethmac_crc32_checker_sink_sink_payload_last_be = ethmac_preamble_checker_source_payload_last_be;
assign ethmac_crc32_checker_sink_sink_payload_error = ethmac_preamble_checker_source_payload_error;
assign ethmac_padding_checker_sink_valid = ethmac_crc32_checker_source_source_valid;
assign ethmac_crc32_checker_source_source_ready = ethmac_padding_checker_sink_ready;
assign ethmac_padding_checker_sink_first = ethmac_crc32_checker_source_source_first;
assign ethmac_padding_checker_sink_last = ethmac_crc32_checker_source_source_last;
assign ethmac_padding_checker_sink_payload_data = ethmac_crc32_checker_source_source_payload_data;
assign ethmac_padding_checker_sink_payload_last_be = ethmac_crc32_checker_source_source_payload_last_be;
assign ethmac_padding_checker_sink_payload_error = ethmac_crc32_checker_source_source_payload_error;
assign ethmac_rx_last_be_sink_valid = ethmac_padding_checker_source_valid;
assign ethmac_padding_checker_source_ready = ethmac_rx_last_be_sink_ready;
assign ethmac_rx_last_be_sink_first = ethmac_padding_checker_source_first;
assign ethmac_rx_last_be_sink_last = ethmac_padding_checker_source_last;
assign ethmac_rx_last_be_sink_payload_data = ethmac_padding_checker_source_payload_data;
assign ethmac_rx_last_be_sink_payload_last_be = ethmac_padding_checker_source_payload_last_be;
assign ethmac_rx_last_be_sink_payload_error = ethmac_padding_checker_source_payload_error;
assign ethmac_rx_converter_sink_valid = ethmac_rx_last_be_source_valid;
assign ethmac_rx_last_be_source_ready = ethmac_rx_converter_sink_ready;
assign ethmac_rx_converter_sink_first = ethmac_rx_last_be_source_first;
assign ethmac_rx_converter_sink_last = ethmac_rx_last_be_source_last;
assign ethmac_rx_converter_sink_payload_data = ethmac_rx_last_be_source_payload_data;
assign ethmac_rx_converter_sink_payload_last_be = ethmac_rx_last_be_source_payload_last_be;
assign ethmac_rx_converter_sink_payload_error = ethmac_rx_last_be_source_payload_error;
assign ethmac_rx_cdc_sink_valid = ethmac_rx_converter_source_valid;
assign ethmac_rx_converter_source_ready = ethmac_rx_cdc_sink_ready;
assign ethmac_rx_cdc_sink_first = ethmac_rx_converter_source_first;
assign ethmac_rx_cdc_sink_last = ethmac_rx_converter_source_last;
assign ethmac_rx_cdc_sink_payload_data = ethmac_rx_converter_source_payload_data;
assign ethmac_rx_cdc_sink_payload_last_be = ethmac_rx_converter_source_payload_last_be;
assign ethmac_rx_cdc_sink_payload_error = ethmac_rx_converter_source_payload_error;
assign ethmac_writer_sink_sink_valid = ethmac_sink_valid;
assign ethmac_sink_ready = ethmac_writer_sink_sink_ready;
assign ethmac_writer_sink_sink_first = ethmac_sink_first;
assign ethmac_writer_sink_sink_last = ethmac_sink_last;
assign ethmac_writer_sink_sink_payload_data = ethmac_sink_payload_data;
assign ethmac_writer_sink_sink_payload_last_be = ethmac_sink_payload_last_be;
assign ethmac_writer_sink_sink_payload_error = ethmac_sink_payload_error;
assign ethmac_source_valid = ethmac_reader_source_source_valid;
assign ethmac_reader_source_source_ready = ethmac_source_ready;
assign ethmac_source_first = ethmac_reader_source_source_first;
assign ethmac_source_last = ethmac_reader_source_source_last;
assign ethmac_source_payload_data = ethmac_reader_source_source_payload_data;
assign ethmac_source_payload_last_be = ethmac_reader_source_source_payload_last_be;
assign ethmac_source_payload_error = ethmac_reader_source_source_payload_error;
always @(*) begin
	ethmac_writer_increment <= 3'd0;
	if (ethmac_writer_sink_sink_payload_last_be[3]) begin
		ethmac_writer_increment <= 1'd1;
	end else begin
		if (ethmac_writer_sink_sink_payload_last_be[2]) begin
			ethmac_writer_increment <= 2'd2;
		end else begin
			if (ethmac_writer_sink_sink_payload_last_be[1]) begin
				ethmac_writer_increment <= 2'd3;
			end else begin
				ethmac_writer_increment <= 3'd4;
			end
		end
	end
end
assign ethmac_writer_fifo_sink_payload_slot = ethmac_writer_slot;
assign ethmac_writer_fifo_sink_payload_length = ethmac_writer_counter;
assign ethmac_writer_fifo_source_ready = ethmac_writer_available_clear;
assign ethmac_writer_available_trigger = ethmac_writer_fifo_source_valid;
assign ethmac_writer_slot_status = ethmac_writer_fifo_source_payload_slot;
assign ethmac_writer_length_status = ethmac_writer_fifo_source_payload_length;
always @(*) begin
	ethmac_writer_memory0_dat_w <= 32'd0;
	ethmac_writer_memory1_adr <= 9'd0;
	ethmac_writer_memory1_we <= 1'd0;
	ethmac_writer_memory0_adr <= 9'd0;
	ethmac_writer_memory1_dat_w <= 32'd0;
	ethmac_writer_memory0_we <= 1'd0;
	case (ethmac_writer_slot)
		1'd0: begin
			ethmac_writer_memory0_adr <= ethmac_writer_counter[31:2];
			ethmac_writer_memory0_dat_w <= ethmac_writer_sink_sink_payload_data;
			if ((ethmac_writer_sink_sink_valid & ethmac_writer_ongoing)) begin
				ethmac_writer_memory0_we <= 4'd15;
			end
		end
		1'd1: begin
			ethmac_writer_memory1_adr <= ethmac_writer_counter[31:2];
			ethmac_writer_memory1_dat_w <= ethmac_writer_sink_sink_payload_data;
			if ((ethmac_writer_sink_sink_valid & ethmac_writer_ongoing)) begin
				ethmac_writer_memory1_we <= 4'd15;
			end
		end
	endcase
end
assign ethmac_writer_status_w = ethmac_writer_available_status;
always @(*) begin
	ethmac_writer_available_clear <= 1'd0;
	if ((ethmac_writer_pending_re & ethmac_writer_pending_r)) begin
		ethmac_writer_available_clear <= 1'd1;
	end
end
assign ethmac_writer_pending_w = ethmac_writer_available_pending;
assign ethmac_writer_irq = (ethmac_writer_pending_w & ethmac_writer_storage);
assign ethmac_writer_available_status = ethmac_writer_available_trigger;
assign ethmac_writer_available_pending = ethmac_writer_available_trigger;
assign ethmac_writer_fifo_syncfifo_din = {ethmac_writer_fifo_fifo_in_last, ethmac_writer_fifo_fifo_in_first, ethmac_writer_fifo_fifo_in_payload_length, ethmac_writer_fifo_fifo_in_payload_slot};
assign {ethmac_writer_fifo_fifo_out_last, ethmac_writer_fifo_fifo_out_first, ethmac_writer_fifo_fifo_out_payload_length, ethmac_writer_fifo_fifo_out_payload_slot} = ethmac_writer_fifo_syncfifo_dout;
assign ethmac_writer_fifo_sink_ready = ethmac_writer_fifo_syncfifo_writable;
assign ethmac_writer_fifo_syncfifo_we = ethmac_writer_fifo_sink_valid;
assign ethmac_writer_fifo_fifo_in_first = ethmac_writer_fifo_sink_first;
assign ethmac_writer_fifo_fifo_in_last = ethmac_writer_fifo_sink_last;
assign ethmac_writer_fifo_fifo_in_payload_slot = ethmac_writer_fifo_sink_payload_slot;
assign ethmac_writer_fifo_fifo_in_payload_length = ethmac_writer_fifo_sink_payload_length;
assign ethmac_writer_fifo_source_valid = ethmac_writer_fifo_syncfifo_readable;
assign ethmac_writer_fifo_source_first = ethmac_writer_fifo_fifo_out_first;
assign ethmac_writer_fifo_source_last = ethmac_writer_fifo_fifo_out_last;
assign ethmac_writer_fifo_source_payload_slot = ethmac_writer_fifo_fifo_out_payload_slot;
assign ethmac_writer_fifo_source_payload_length = ethmac_writer_fifo_fifo_out_payload_length;
assign ethmac_writer_fifo_syncfifo_re = ethmac_writer_fifo_source_ready;
always @(*) begin
	ethmac_writer_fifo_wrport_adr <= 1'd0;
	if (ethmac_writer_fifo_replace) begin
		ethmac_writer_fifo_wrport_adr <= (ethmac_writer_fifo_produce - 1'd1);
	end else begin
		ethmac_writer_fifo_wrport_adr <= ethmac_writer_fifo_produce;
	end
end
assign ethmac_writer_fifo_wrport_dat_w = ethmac_writer_fifo_syncfifo_din;
assign ethmac_writer_fifo_wrport_we = (ethmac_writer_fifo_syncfifo_we & (ethmac_writer_fifo_syncfifo_writable | ethmac_writer_fifo_replace));
assign ethmac_writer_fifo_do_read = (ethmac_writer_fifo_syncfifo_readable & ethmac_writer_fifo_syncfifo_re);
assign ethmac_writer_fifo_rdport_adr = ethmac_writer_fifo_consume;
assign ethmac_writer_fifo_syncfifo_dout = ethmac_writer_fifo_rdport_dat_r;
assign ethmac_writer_fifo_syncfifo_writable = (ethmac_writer_fifo_level != 2'd2);
assign ethmac_writer_fifo_syncfifo_readable = (ethmac_writer_fifo_level != 1'd0);
always @(*) begin
	ethmac_writer_counter_reset <= 1'd0;
	ethmac_writer_counter_ce <= 1'd0;
	liteethmacsramwriter_next_state <= 3'd0;
	ethmac_writer_errors_status_liteethmac_next_value <= 32'd0;
	ethmac_writer_slot_ce <= 1'd0;
	ethmac_writer_errors_status_liteethmac_next_value_ce <= 1'd0;
	ethmac_writer_ongoing <= 1'd0;
	ethmac_writer_fifo_sink_valid <= 1'd0;
	liteethmacsramwriter_next_state <= liteethmacsramwriter_state;
	case (liteethmacsramwriter_state)
		1'd1: begin
			if (ethmac_writer_sink_sink_valid) begin
				if ((ethmac_writer_counter == 11'd1530)) begin
					liteethmacsramwriter_next_state <= 2'd3;
				end else begin
					ethmac_writer_counter_ce <= 1'd1;
					ethmac_writer_ongoing <= 1'd1;
				end
				if (ethmac_writer_sink_sink_last) begin
					if (((ethmac_writer_sink_sink_payload_error & ethmac_writer_sink_sink_payload_last_be) != 1'd0)) begin
						liteethmacsramwriter_next_state <= 2'd2;
					end else begin
						liteethmacsramwriter_next_state <= 3'd4;
					end
				end
			end
		end
		2'd2: begin
			ethmac_writer_counter_reset <= 1'd1;
			liteethmacsramwriter_next_state <= 1'd0;
		end
		2'd3: begin
			if ((ethmac_writer_sink_sink_valid & ethmac_writer_sink_sink_last)) begin
				liteethmacsramwriter_next_state <= 3'd4;
			end
		end
		3'd4: begin
			ethmac_writer_counter_reset <= 1'd1;
			ethmac_writer_slot_ce <= 1'd1;
			ethmac_writer_fifo_sink_valid <= 1'd1;
			liteethmacsramwriter_next_state <= 1'd0;
		end
		default: begin
			if (ethmac_writer_sink_sink_valid) begin
				if (ethmac_writer_fifo_sink_ready) begin
					ethmac_writer_ongoing <= 1'd1;
					ethmac_writer_counter_ce <= 1'd1;
					liteethmacsramwriter_next_state <= 1'd1;
				end else begin
					ethmac_writer_errors_status_liteethmac_next_value <= (ethmac_writer_errors_status + 1'd1);
					ethmac_writer_errors_status_liteethmac_next_value_ce <= 1'd1;
					liteethmacsramwriter_next_state <= 2'd3;
				end
			end
		end
	endcase
end
assign ethmac_reader_fifo_sink_valid = ethmac_reader_start_re;
assign ethmac_reader_fifo_sink_payload_slot = ethmac_reader_slot_storage;
assign ethmac_reader_fifo_sink_payload_length = ethmac_reader_length_storage;
assign ethmac_reader_ready_status = ethmac_reader_fifo_sink_ready;
assign ethmac_reader_level_status = ethmac_reader_fifo_level;
always @(*) begin
	ethmac_reader_source_source_payload_last_be <= 4'd0;
	if (ethmac_reader_last) begin
		if ((ethmac_reader_fifo_source_payload_length[1:0] == 2'd3)) begin
			ethmac_reader_source_source_payload_last_be <= 2'd2;
		end else begin
			if ((ethmac_reader_fifo_source_payload_length[1:0] == 2'd2)) begin
				ethmac_reader_source_source_payload_last_be <= 3'd4;
			end else begin
				if ((ethmac_reader_fifo_source_payload_length[1:0] == 1'd1)) begin
					ethmac_reader_source_source_payload_last_be <= 4'd8;
				end else begin
					ethmac_reader_source_source_payload_last_be <= 1'd1;
				end
			end
		end
	end
end
assign ethmac_reader_last = ((ethmac_reader_counter + 3'd4) >= ethmac_reader_fifo_source_payload_length);
assign ethmac_reader_memory0_adr = ethmac_reader_counter[10:2];
assign ethmac_reader_memory1_adr = ethmac_reader_counter[10:2];
always @(*) begin
	ethmac_reader_source_source_payload_data <= 32'd0;
	case (ethmac_reader_fifo_source_payload_slot)
		1'd0: begin
			ethmac_reader_source_source_payload_data <= ethmac_reader_memory0_dat_r;
		end
		1'd1: begin
			ethmac_reader_source_source_payload_data <= ethmac_reader_memory1_dat_r;
		end
	endcase
end
assign ethmac_reader_eventmanager_status_w = ethmac_reader_done_status;
always @(*) begin
	ethmac_reader_done_clear <= 1'd0;
	if ((ethmac_reader_eventmanager_pending_re & ethmac_reader_eventmanager_pending_r)) begin
		ethmac_reader_done_clear <= 1'd1;
	end
end
assign ethmac_reader_eventmanager_pending_w = ethmac_reader_done_pending;
assign ethmac_reader_irq = (ethmac_reader_eventmanager_pending_w & ethmac_reader_eventmanager_storage);
assign ethmac_reader_done_status = 1'd0;
assign ethmac_reader_fifo_syncfifo_din = {ethmac_reader_fifo_fifo_in_last, ethmac_reader_fifo_fifo_in_first, ethmac_reader_fifo_fifo_in_payload_length, ethmac_reader_fifo_fifo_in_payload_slot};
assign {ethmac_reader_fifo_fifo_out_last, ethmac_reader_fifo_fifo_out_first, ethmac_reader_fifo_fifo_out_payload_length, ethmac_reader_fifo_fifo_out_payload_slot} = ethmac_reader_fifo_syncfifo_dout;
assign ethmac_reader_fifo_sink_ready = ethmac_reader_fifo_syncfifo_writable;
assign ethmac_reader_fifo_syncfifo_we = ethmac_reader_fifo_sink_valid;
assign ethmac_reader_fifo_fifo_in_first = ethmac_reader_fifo_sink_first;
assign ethmac_reader_fifo_fifo_in_last = ethmac_reader_fifo_sink_last;
assign ethmac_reader_fifo_fifo_in_payload_slot = ethmac_reader_fifo_sink_payload_slot;
assign ethmac_reader_fifo_fifo_in_payload_length = ethmac_reader_fifo_sink_payload_length;
assign ethmac_reader_fifo_source_valid = ethmac_reader_fifo_syncfifo_readable;
assign ethmac_reader_fifo_source_first = ethmac_reader_fifo_fifo_out_first;
assign ethmac_reader_fifo_source_last = ethmac_reader_fifo_fifo_out_last;
assign ethmac_reader_fifo_source_payload_slot = ethmac_reader_fifo_fifo_out_payload_slot;
assign ethmac_reader_fifo_source_payload_length = ethmac_reader_fifo_fifo_out_payload_length;
assign ethmac_reader_fifo_syncfifo_re = ethmac_reader_fifo_source_ready;
always @(*) begin
	ethmac_reader_fifo_wrport_adr <= 1'd0;
	if (ethmac_reader_fifo_replace) begin
		ethmac_reader_fifo_wrport_adr <= (ethmac_reader_fifo_produce - 1'd1);
	end else begin
		ethmac_reader_fifo_wrport_adr <= ethmac_reader_fifo_produce;
	end
end
assign ethmac_reader_fifo_wrport_dat_w = ethmac_reader_fifo_syncfifo_din;
assign ethmac_reader_fifo_wrport_we = (ethmac_reader_fifo_syncfifo_we & (ethmac_reader_fifo_syncfifo_writable | ethmac_reader_fifo_replace));
assign ethmac_reader_fifo_do_read = (ethmac_reader_fifo_syncfifo_readable & ethmac_reader_fifo_syncfifo_re);
assign ethmac_reader_fifo_rdport_adr = ethmac_reader_fifo_consume;
assign ethmac_reader_fifo_syncfifo_dout = ethmac_reader_fifo_rdport_dat_r;
assign ethmac_reader_fifo_syncfifo_writable = (ethmac_reader_fifo_level != 2'd2);
assign ethmac_reader_fifo_syncfifo_readable = (ethmac_reader_fifo_level != 1'd0);
always @(*) begin
	liteethmacsramreader_next_state <= 2'd0;
	ethmac_reader_done_trigger <= 1'd0;
	ethmac_reader_source_source_valid <= 1'd0;
	ethmac_reader_counter_reset <= 1'd0;
	ethmac_reader_counter_ce <= 1'd0;
	ethmac_reader_fifo_source_ready <= 1'd0;
	ethmac_reader_source_source_last <= 1'd0;
	liteethmacsramreader_next_state <= liteethmacsramreader_state;
	case (liteethmacsramreader_state)
		1'd1: begin
			if ((~ethmac_reader_last_d)) begin
				liteethmacsramreader_next_state <= 2'd2;
			end else begin
				liteethmacsramreader_next_state <= 2'd3;
			end
		end
		2'd2: begin
			ethmac_reader_source_source_valid <= 1'd1;
			ethmac_reader_source_source_last <= ethmac_reader_last;
			if (ethmac_reader_source_source_ready) begin
				ethmac_reader_counter_ce <= (~ethmac_reader_last);
				liteethmacsramreader_next_state <= 1'd1;
			end
		end
		2'd3: begin
			ethmac_reader_fifo_source_ready <= 1'd1;
			ethmac_reader_done_trigger <= 1'd1;
			liteethmacsramreader_next_state <= 1'd0;
		end
		default: begin
			ethmac_reader_counter_reset <= 1'd1;
			if (ethmac_reader_fifo_source_valid) begin
				liteethmacsramreader_next_state <= 1'd1;
			end
		end
	endcase
end
assign ethmac_ev_irq = (ethmac_writer_irq | ethmac_reader_irq);
assign ethmac_sram0_adr0 = ethmac_sram0_bus_adr0[8:0];
assign ethmac_sram0_bus_dat_r0 = ethmac_sram0_dat_r0;
assign ethmac_sram1_adr0 = ethmac_sram1_bus_adr0[8:0];
assign ethmac_sram1_bus_dat_r0 = ethmac_sram1_dat_r0;
always @(*) begin
	ethmac_sram0_we <= 4'd0;
	ethmac_sram0_we[0] <= (((ethmac_sram0_bus_cyc1 & ethmac_sram0_bus_stb1) & ethmac_sram0_bus_we1) & ethmac_sram0_bus_sel1[0]);
	ethmac_sram0_we[1] <= (((ethmac_sram0_bus_cyc1 & ethmac_sram0_bus_stb1) & ethmac_sram0_bus_we1) & ethmac_sram0_bus_sel1[1]);
	ethmac_sram0_we[2] <= (((ethmac_sram0_bus_cyc1 & ethmac_sram0_bus_stb1) & ethmac_sram0_bus_we1) & ethmac_sram0_bus_sel1[2]);
	ethmac_sram0_we[3] <= (((ethmac_sram0_bus_cyc1 & ethmac_sram0_bus_stb1) & ethmac_sram0_bus_we1) & ethmac_sram0_bus_sel1[3]);
end
assign ethmac_sram0_adr1 = ethmac_sram0_bus_adr1[8:0];
assign ethmac_sram0_bus_dat_r1 = ethmac_sram0_dat_r1;
assign ethmac_sram0_dat_w = ethmac_sram0_bus_dat_w1;
always @(*) begin
	ethmac_sram1_we <= 4'd0;
	ethmac_sram1_we[0] <= (((ethmac_sram1_bus_cyc1 & ethmac_sram1_bus_stb1) & ethmac_sram1_bus_we1) & ethmac_sram1_bus_sel1[0]);
	ethmac_sram1_we[1] <= (((ethmac_sram1_bus_cyc1 & ethmac_sram1_bus_stb1) & ethmac_sram1_bus_we1) & ethmac_sram1_bus_sel1[1]);
	ethmac_sram1_we[2] <= (((ethmac_sram1_bus_cyc1 & ethmac_sram1_bus_stb1) & ethmac_sram1_bus_we1) & ethmac_sram1_bus_sel1[2]);
	ethmac_sram1_we[3] <= (((ethmac_sram1_bus_cyc1 & ethmac_sram1_bus_stb1) & ethmac_sram1_bus_we1) & ethmac_sram1_bus_sel1[3]);
end
assign ethmac_sram1_adr1 = ethmac_sram1_bus_adr1[8:0];
assign ethmac_sram1_bus_dat_r1 = ethmac_sram1_dat_r1;
assign ethmac_sram1_dat_w = ethmac_sram1_bus_dat_w1;
always @(*) begin
	ethmac_slave_sel <= 4'd0;
	ethmac_slave_sel[0] <= (ethmac_bus_adr[10:9] == 1'd0);
	ethmac_slave_sel[1] <= (ethmac_bus_adr[10:9] == 1'd1);
	ethmac_slave_sel[2] <= (ethmac_bus_adr[10:9] == 2'd2);
	ethmac_slave_sel[3] <= (ethmac_bus_adr[10:9] == 2'd3);
end
assign ethmac_sram0_bus_adr0 = ethmac_bus_adr;
assign ethmac_sram0_bus_dat_w0 = ethmac_bus_dat_w;
assign ethmac_sram0_bus_sel0 = ethmac_bus_sel;
assign ethmac_sram0_bus_stb0 = ethmac_bus_stb;
assign ethmac_sram0_bus_we0 = ethmac_bus_we;
assign ethmac_sram0_bus_cti0 = ethmac_bus_cti;
assign ethmac_sram0_bus_bte0 = ethmac_bus_bte;
assign ethmac_sram1_bus_adr0 = ethmac_bus_adr;
assign ethmac_sram1_bus_dat_w0 = ethmac_bus_dat_w;
assign ethmac_sram1_bus_sel0 = ethmac_bus_sel;
assign ethmac_sram1_bus_stb0 = ethmac_bus_stb;
assign ethmac_sram1_bus_we0 = ethmac_bus_we;
assign ethmac_sram1_bus_cti0 = ethmac_bus_cti;
assign ethmac_sram1_bus_bte0 = ethmac_bus_bte;
assign ethmac_sram0_bus_adr1 = ethmac_bus_adr;
assign ethmac_sram0_bus_dat_w1 = ethmac_bus_dat_w;
assign ethmac_sram0_bus_sel1 = ethmac_bus_sel;
assign ethmac_sram0_bus_stb1 = ethmac_bus_stb;
assign ethmac_sram0_bus_we1 = ethmac_bus_we;
assign ethmac_sram0_bus_cti1 = ethmac_bus_cti;
assign ethmac_sram0_bus_bte1 = ethmac_bus_bte;
assign ethmac_sram1_bus_adr1 = ethmac_bus_adr;
assign ethmac_sram1_bus_dat_w1 = ethmac_bus_dat_w;
assign ethmac_sram1_bus_sel1 = ethmac_bus_sel;
assign ethmac_sram1_bus_stb1 = ethmac_bus_stb;
assign ethmac_sram1_bus_we1 = ethmac_bus_we;
assign ethmac_sram1_bus_cti1 = ethmac_bus_cti;
assign ethmac_sram1_bus_bte1 = ethmac_bus_bte;
assign ethmac_sram0_bus_cyc0 = (ethmac_bus_cyc & ethmac_slave_sel[0]);
assign ethmac_sram1_bus_cyc0 = (ethmac_bus_cyc & ethmac_slave_sel[1]);
assign ethmac_sram0_bus_cyc1 = (ethmac_bus_cyc & ethmac_slave_sel[2]);
assign ethmac_sram1_bus_cyc1 = (ethmac_bus_cyc & ethmac_slave_sel[3]);
assign ethmac_bus_ack = (((ethmac_sram0_bus_ack0 | ethmac_sram1_bus_ack0) | ethmac_sram0_bus_ack1) | ethmac_sram1_bus_ack1);
assign ethmac_bus_err = (((ethmac_sram0_bus_err0 | ethmac_sram1_bus_err0) | ethmac_sram0_bus_err1) | ethmac_sram1_bus_err1);
assign ethmac_bus_dat_r = (((({32{ethmac_slave_sel_r[0]}} & ethmac_sram0_bus_dat_r0) | ({32{ethmac_slave_sel_r[1]}} & ethmac_sram1_bus_dat_r0)) | ({32{ethmac_slave_sel_r[2]}} & ethmac_sram0_bus_dat_r1)) | ({32{ethmac_slave_sel_r[3]}} & ethmac_sram1_bus_dat_r1));
assign charsync0_raw_data = s7datacapture0_d;
assign wer0_data = charsync0_data;
assign decoding0_valid_i = charsync0_synced;
assign decoding0_input = charsync0_data;
assign charsync1_raw_data = s7datacapture1_d;
assign wer1_data = charsync1_data;
assign decoding1_valid_i = charsync1_synced;
assign decoding1_input = charsync1_data;
assign charsync2_raw_data = s7datacapture2_d;
assign wer2_data = charsync2_data;
assign decoding2_valid_i = charsync2_synced;
assign decoding2_input = charsync2_data;
assign chansync_valid_i = ((decoding0_valid_o & decoding1_valid_o) & decoding2_valid_o);
assign chansync_data_in0_d = decoding0_output_d;
assign chansync_data_in0_c = decoding0_output_c;
assign chansync_data_in0_de = decoding0_output_de;
assign chansync_data_in1_d = decoding1_output_d;
assign chansync_data_in1_c = decoding1_output_c;
assign chansync_data_in1_de = decoding1_output_de;
assign chansync_data_in2_d = decoding2_output_d;
assign chansync_data_in2_c = decoding2_output_c;
assign chansync_data_in2_de = decoding2_output_de;
assign syncpol_valid_i = chansync_chan_synced;
assign syncpol_data_in0_d = chansync_data_out0_d;
assign syncpol_data_in0_c = chansync_data_out0_c;
assign syncpol_data_in0_de = chansync_data_out0_de;
assign syncpol_data_in1_d = chansync_data_out1_d;
assign syncpol_data_in1_c = chansync_data_out1_c;
assign syncpol_data_in1_de = chansync_data_out1_de;
assign syncpol_data_in2_d = chansync_data_out2_d;
assign syncpol_data_in2_c = chansync_data_out2_c;
assign syncpol_data_in2_de = chansync_data_out2_de;
assign resdetection_valid_i = syncpol_valid_o;
assign resdetection_de = syncpol_de;
assign resdetection_vsync = syncpol_vsync;
assign frame_valid_i = syncpol_valid_o;
assign frame_de = syncpol_de;
assign frame_vsync = syncpol_vsync;
assign frame_r = syncpol_r;
assign frame_g = syncpol_g;
assign frame_b = syncpol_b;
assign dma_frame_valid = frame_frame_valid;
assign frame_frame_ready = dma_frame_ready;
assign dma_frame_first = frame_frame_first;
assign dma_frame_last = frame_frame_last;
assign dma_frame_payload_sof = frame_frame_payload_sof;
assign dma_frame_payload_pixels = frame_frame_payload_pixels;
assign edid_status = 1'd1;
assign hdmi_in_hpd_en = edid_storage;
assign edid_sda_o = (~edid_sda_drv_reg);
assign edid_scl_rising = (edid_scl_i & (~edid_scl_r));
assign edid_sda_rising = (edid_sda_i & (~edid_sda_r));
assign edid_sda_falling = ((~edid_sda_i) & edid_sda_r);
assign edid_start = (edid_scl_i & edid_sda_falling);
assign edid_adr = edid_offset_counter;
always @(*) begin
	edid_sda_drv <= 1'd0;
	if (edid_zero_drv) begin
		edid_sda_drv <= 1'd1;
	end else begin
		if (edid_data_drv) begin
			edid_sda_drv <= (~edid_data_bit);
		end
	end
end
always @(*) begin
	edid_update_is_read <= 1'd0;
	edid_zero_drv <= 1'd0;
	edid_oc_load <= 1'd0;
	edid_oc_inc <= 1'd0;
	edid_data_drv_en <= 1'd0;
	edid_data_drv_stop <= 1'd0;
	edid_next_state <= 4'd0;
	edid_next_state <= edid_state;
	case (edid_state)
		1'd1: begin
			if ((edid_counter == 4'd8)) begin
				if ((edid_din[7:1] == 7'd80)) begin
					edid_update_is_read <= 1'd1;
					edid_next_state <= 2'd2;
				end else begin
					edid_next_state <= 1'd0;
				end
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		2'd2: begin
			if ((~edid_scl_i)) begin
				edid_next_state <= 2'd3;
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		2'd3: begin
			edid_zero_drv <= 1'd1;
			if (edid_scl_i) begin
				edid_next_state <= 3'd4;
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		3'd4: begin
			edid_zero_drv <= 1'd1;
			if ((~edid_scl_i)) begin
				if (edid_is_read) begin
					edid_next_state <= 4'd9;
				end else begin
					edid_next_state <= 3'd5;
				end
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		3'd5: begin
			if ((edid_counter == 4'd8)) begin
				edid_oc_load <= 1'd1;
				edid_next_state <= 3'd6;
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		3'd6: begin
			if ((~edid_scl_i)) begin
				edid_next_state <= 3'd7;
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		3'd7: begin
			edid_zero_drv <= 1'd1;
			if (edid_scl_i) begin
				edid_next_state <= 4'd8;
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		4'd8: begin
			edid_zero_drv <= 1'd1;
			if ((~edid_scl_i)) begin
				edid_next_state <= 1'd1;
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		4'd9: begin
			if ((~edid_scl_i)) begin
				if ((edid_counter == 4'd8)) begin
					edid_data_drv_stop <= 1'd1;
					edid_next_state <= 4'd10;
				end else begin
					edid_data_drv_en <= 1'd1;
				end
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		4'd10: begin
			if (edid_scl_rising) begin
				edid_oc_inc <= 1'd1;
				if (edid_sda_i) begin
					edid_next_state <= 1'd0;
				end else begin
					edid_next_state <= 4'd9;
				end
			end
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
		default: begin
			if (edid_start) begin
				edid_next_state <= 1'd1;
			end
			if ((~edid_storage)) begin
				edid_next_state <= 1'd0;
			end
		end
	endcase
end
assign locked_status = locked;
assign s7datacapture0_serdes_m_d = s7datacapture0_serdes_m_q;
assign s7datacapture0_serdes_s_d = s7datacapture0_serdes_s_q;
assign s7datacapture0_gearbox_i = s7datacapture0_serdes_m_d;
assign s7datacapture0_d = s7datacapture0_gearbox_o;
assign s7datacapture0_mdata = s7datacapture0_serdes_m_d;
assign s7datacapture0_sdata = (~s7datacapture0_serdes_s_d);
assign s7datacapture0_too_late = (s7datacapture0_lateness == 8'd255);
assign s7datacapture0_too_early = (s7datacapture0_lateness == 1'd0);
assign s7datacapture0_delay_rst = s7datacapture0_do_delay_rst_o;
assign s7datacapture0_delay_master_inc = s7datacapture0_do_delay_master_inc_o;
assign s7datacapture0_delay_master_ce = (s7datacapture0_do_delay_master_inc_o | s7datacapture0_do_delay_master_dec_o);
assign s7datacapture0_delay_slave_inc = s7datacapture0_do_delay_slave_inc_o;
assign s7datacapture0_delay_slave_ce = (s7datacapture0_do_delay_slave_inc_o | s7datacapture0_do_delay_slave_dec_o);
assign s7datacapture0_do_delay_rst_i = (s7datacapture0_dly_ctl_re & s7datacapture0_dly_ctl_r[0]);
assign s7datacapture0_do_delay_master_inc_i = (s7datacapture0_dly_ctl_re & s7datacapture0_dly_ctl_r[1]);
assign s7datacapture0_do_delay_master_dec_i = (s7datacapture0_dly_ctl_re & s7datacapture0_dly_ctl_r[2]);
assign s7datacapture0_do_delay_slave_inc_i = (s7datacapture0_dly_ctl_re & s7datacapture0_dly_ctl_r[3]);
assign s7datacapture0_do_delay_slave_dec_i = (s7datacapture0_dly_ctl_re & s7datacapture0_dly_ctl_r[4]);
assign s7datacapture0_reset_lateness = s7datacapture0_do_reset_lateness_o;
assign s7datacapture0_do_reset_lateness_i = s7datacapture0_phase_reset_re;
assign s7datacapture0_gearbox_rst = (pix1p25x_rst | hdmi_in0_pix_rst);
assign data0_cap_write_clk = pix1p25x_clk;
assign data0_cap_read_clk = hdmi_in0_pix_clk;
assign data0_cap_write_rst = s7datacapture0_gearbox_rst;
assign data0_cap_read_rst = s7datacapture0_gearbox_rst;
assign s7datacapture0_transition = (s7datacapture0_mdata_d != s7datacapture0_mdata);
assign s7datacapture0_inc = (s7datacapture0_transition & (s7datacapture0_mdata == s7datacapture0_sdata));
assign s7datacapture0_dec = (s7datacapture0_transition & (s7datacapture0_mdata != s7datacapture0_sdata));
assign s7datacapture0_do_delay_rst_o = (s7datacapture0_do_delay_rst_toggle_o ^ s7datacapture0_do_delay_rst_toggle_o_r);
assign s7datacapture0_do_delay_master_inc_o = (s7datacapture0_do_delay_master_inc_toggle_o ^ s7datacapture0_do_delay_master_inc_toggle_o_r);
assign s7datacapture0_do_delay_master_dec_o = (s7datacapture0_do_delay_master_dec_toggle_o ^ s7datacapture0_do_delay_master_dec_toggle_o_r);
assign s7datacapture0_do_delay_slave_inc_o = (s7datacapture0_do_delay_slave_inc_toggle_o ^ s7datacapture0_do_delay_slave_inc_toggle_o_r);
assign s7datacapture0_do_delay_slave_dec_o = (s7datacapture0_do_delay_slave_dec_toggle_o ^ s7datacapture0_do_delay_slave_dec_toggle_o_r);
assign s7datacapture0_do_reset_lateness_o = (s7datacapture0_do_reset_lateness_toggle_o ^ s7datacapture0_do_reset_lateness_toggle_o_r);
assign charsync0_raw = {charsync0_raw_data, charsync0_raw_data1};
always @(*) begin
	wer0_transitions <= 8'd0;
	wer0_transitions[0] <= (wer0_data_r[0] ^ wer0_data_r[1]);
	wer0_transitions[1] <= (wer0_data_r[1] ^ wer0_data_r[2]);
	wer0_transitions[2] <= (wer0_data_r[2] ^ wer0_data_r[3]);
	wer0_transitions[3] <= (wer0_data_r[3] ^ wer0_data_r[4]);
	wer0_transitions[4] <= (wer0_data_r[4] ^ wer0_data_r[5]);
	wer0_transitions[5] <= (wer0_data_r[5] ^ wer0_data_r[6]);
	wer0_transitions[6] <= (wer0_data_r[6] ^ wer0_data_r[7]);
	wer0_transitions[7] <= (wer0_data_r[7] ^ wer0_data_r[8]);
end
assign wer0_i = wer0_wer_counter_r_updated;
assign wer0_o = (wer0_toggle_o ^ wer0_toggle_o_r);
assign s7datacapture1_serdes_m_d = s7datacapture1_serdes_m_q;
assign s7datacapture1_serdes_s_d = s7datacapture1_serdes_s_q;
assign s7datacapture1_gearbox_i = s7datacapture1_serdes_m_d;
assign s7datacapture1_d = s7datacapture1_gearbox_o;
assign s7datacapture1_mdata = s7datacapture1_serdes_m_d;
assign s7datacapture1_sdata = (~s7datacapture1_serdes_s_d);
assign s7datacapture1_too_late = (s7datacapture1_lateness == 8'd255);
assign s7datacapture1_too_early = (s7datacapture1_lateness == 1'd0);
assign s7datacapture1_delay_rst = s7datacapture1_do_delay_rst_o;
assign s7datacapture1_delay_master_inc = s7datacapture1_do_delay_master_inc_o;
assign s7datacapture1_delay_master_ce = (s7datacapture1_do_delay_master_inc_o | s7datacapture1_do_delay_master_dec_o);
assign s7datacapture1_delay_slave_inc = s7datacapture1_do_delay_slave_inc_o;
assign s7datacapture1_delay_slave_ce = (s7datacapture1_do_delay_slave_inc_o | s7datacapture1_do_delay_slave_dec_o);
assign s7datacapture1_do_delay_rst_i = (s7datacapture1_dly_ctl_re & s7datacapture1_dly_ctl_r[0]);
assign s7datacapture1_do_delay_master_inc_i = (s7datacapture1_dly_ctl_re & s7datacapture1_dly_ctl_r[1]);
assign s7datacapture1_do_delay_master_dec_i = (s7datacapture1_dly_ctl_re & s7datacapture1_dly_ctl_r[2]);
assign s7datacapture1_do_delay_slave_inc_i = (s7datacapture1_dly_ctl_re & s7datacapture1_dly_ctl_r[3]);
assign s7datacapture1_do_delay_slave_dec_i = (s7datacapture1_dly_ctl_re & s7datacapture1_dly_ctl_r[4]);
assign s7datacapture1_reset_lateness = s7datacapture1_do_reset_lateness_o;
assign s7datacapture1_do_reset_lateness_i = s7datacapture1_phase_reset_re;
assign s7datacapture1_gearbox_rst = (pix1p25x_rst | hdmi_in0_pix_rst);
assign data1_cap_write_clk = pix1p25x_clk;
assign data1_cap_read_clk = hdmi_in0_pix_clk;
assign data1_cap_write_rst = s7datacapture1_gearbox_rst;
assign data1_cap_read_rst = s7datacapture1_gearbox_rst;
assign s7datacapture1_transition = (s7datacapture1_mdata_d != s7datacapture1_mdata);
assign s7datacapture1_inc = (s7datacapture1_transition & (s7datacapture1_mdata == s7datacapture1_sdata));
assign s7datacapture1_dec = (s7datacapture1_transition & (s7datacapture1_mdata != s7datacapture1_sdata));
assign s7datacapture1_do_delay_rst_o = (s7datacapture1_do_delay_rst_toggle_o ^ s7datacapture1_do_delay_rst_toggle_o_r);
assign s7datacapture1_do_delay_master_inc_o = (s7datacapture1_do_delay_master_inc_toggle_o ^ s7datacapture1_do_delay_master_inc_toggle_o_r);
assign s7datacapture1_do_delay_master_dec_o = (s7datacapture1_do_delay_master_dec_toggle_o ^ s7datacapture1_do_delay_master_dec_toggle_o_r);
assign s7datacapture1_do_delay_slave_inc_o = (s7datacapture1_do_delay_slave_inc_toggle_o ^ s7datacapture1_do_delay_slave_inc_toggle_o_r);
assign s7datacapture1_do_delay_slave_dec_o = (s7datacapture1_do_delay_slave_dec_toggle_o ^ s7datacapture1_do_delay_slave_dec_toggle_o_r);
assign s7datacapture1_do_reset_lateness_o = (s7datacapture1_do_reset_lateness_toggle_o ^ s7datacapture1_do_reset_lateness_toggle_o_r);
assign charsync1_raw = {charsync1_raw_data, charsync1_raw_data1};
always @(*) begin
	wer1_transitions <= 8'd0;
	wer1_transitions[0] <= (wer1_data_r[0] ^ wer1_data_r[1]);
	wer1_transitions[1] <= (wer1_data_r[1] ^ wer1_data_r[2]);
	wer1_transitions[2] <= (wer1_data_r[2] ^ wer1_data_r[3]);
	wer1_transitions[3] <= (wer1_data_r[3] ^ wer1_data_r[4]);
	wer1_transitions[4] <= (wer1_data_r[4] ^ wer1_data_r[5]);
	wer1_transitions[5] <= (wer1_data_r[5] ^ wer1_data_r[6]);
	wer1_transitions[6] <= (wer1_data_r[6] ^ wer1_data_r[7]);
	wer1_transitions[7] <= (wer1_data_r[7] ^ wer1_data_r[8]);
end
assign wer1_i = wer1_wer_counter_r_updated;
assign wer1_o = (wer1_toggle_o ^ wer1_toggle_o_r);
assign s7datacapture2_serdes_m_d = s7datacapture2_serdes_m_q;
assign s7datacapture2_serdes_s_d = s7datacapture2_serdes_s_q;
assign s7datacapture2_gearbox_i = s7datacapture2_serdes_m_d;
assign s7datacapture2_d = s7datacapture2_gearbox_o;
assign s7datacapture2_mdata = s7datacapture2_serdes_m_d;
assign s7datacapture2_sdata = (~s7datacapture2_serdes_s_d);
assign s7datacapture2_too_late = (s7datacapture2_lateness == 8'd255);
assign s7datacapture2_too_early = (s7datacapture2_lateness == 1'd0);
assign s7datacapture2_delay_rst = s7datacapture2_do_delay_rst_o;
assign s7datacapture2_delay_master_inc = s7datacapture2_do_delay_master_inc_o;
assign s7datacapture2_delay_master_ce = (s7datacapture2_do_delay_master_inc_o | s7datacapture2_do_delay_master_dec_o);
assign s7datacapture2_delay_slave_inc = s7datacapture2_do_delay_slave_inc_o;
assign s7datacapture2_delay_slave_ce = (s7datacapture2_do_delay_slave_inc_o | s7datacapture2_do_delay_slave_dec_o);
assign s7datacapture2_do_delay_rst_i = (s7datacapture2_dly_ctl_re & s7datacapture2_dly_ctl_r[0]);
assign s7datacapture2_do_delay_master_inc_i = (s7datacapture2_dly_ctl_re & s7datacapture2_dly_ctl_r[1]);
assign s7datacapture2_do_delay_master_dec_i = (s7datacapture2_dly_ctl_re & s7datacapture2_dly_ctl_r[2]);
assign s7datacapture2_do_delay_slave_inc_i = (s7datacapture2_dly_ctl_re & s7datacapture2_dly_ctl_r[3]);
assign s7datacapture2_do_delay_slave_dec_i = (s7datacapture2_dly_ctl_re & s7datacapture2_dly_ctl_r[4]);
assign s7datacapture2_reset_lateness = s7datacapture2_do_reset_lateness_o;
assign s7datacapture2_do_reset_lateness_i = s7datacapture2_phase_reset_re;
assign s7datacapture2_gearbox_rst = (pix1p25x_rst | hdmi_in0_pix_rst);
assign data2_cap_write_clk = pix1p25x_clk;
assign data2_cap_read_clk = hdmi_in0_pix_clk;
assign data2_cap_write_rst = s7datacapture2_gearbox_rst;
assign data2_cap_read_rst = s7datacapture2_gearbox_rst;
assign s7datacapture2_transition = (s7datacapture2_mdata_d != s7datacapture2_mdata);
assign s7datacapture2_inc = (s7datacapture2_transition & (s7datacapture2_mdata == s7datacapture2_sdata));
assign s7datacapture2_dec = (s7datacapture2_transition & (s7datacapture2_mdata != s7datacapture2_sdata));
assign s7datacapture2_do_delay_rst_o = (s7datacapture2_do_delay_rst_toggle_o ^ s7datacapture2_do_delay_rst_toggle_o_r);
assign s7datacapture2_do_delay_master_inc_o = (s7datacapture2_do_delay_master_inc_toggle_o ^ s7datacapture2_do_delay_master_inc_toggle_o_r);
assign s7datacapture2_do_delay_master_dec_o = (s7datacapture2_do_delay_master_dec_toggle_o ^ s7datacapture2_do_delay_master_dec_toggle_o_r);
assign s7datacapture2_do_delay_slave_inc_o = (s7datacapture2_do_delay_slave_inc_toggle_o ^ s7datacapture2_do_delay_slave_inc_toggle_o_r);
assign s7datacapture2_do_delay_slave_dec_o = (s7datacapture2_do_delay_slave_dec_toggle_o ^ s7datacapture2_do_delay_slave_dec_toggle_o_r);
assign s7datacapture2_do_reset_lateness_o = (s7datacapture2_do_reset_lateness_toggle_o ^ s7datacapture2_do_reset_lateness_toggle_o_r);
assign charsync2_raw = {charsync2_raw_data, charsync2_raw_data1};
always @(*) begin
	wer2_transitions <= 8'd0;
	wer2_transitions[0] <= (wer2_data_r[0] ^ wer2_data_r[1]);
	wer2_transitions[1] <= (wer2_data_r[1] ^ wer2_data_r[2]);
	wer2_transitions[2] <= (wer2_data_r[2] ^ wer2_data_r[3]);
	wer2_transitions[3] <= (wer2_data_r[3] ^ wer2_data_r[4]);
	wer2_transitions[4] <= (wer2_data_r[4] ^ wer2_data_r[5]);
	wer2_transitions[5] <= (wer2_data_r[5] ^ wer2_data_r[6]);
	wer2_transitions[6] <= (wer2_data_r[6] ^ wer2_data_r[7]);
	wer2_transitions[7] <= (wer2_data_r[7] ^ wer2_data_r[8]);
end
assign wer2_i = wer2_wer_counter_r_updated;
assign wer2_o = (wer2_toggle_o ^ wer2_toggle_o_r);
assign chansync_syncbuffer0_din = {chansync_data_in0_de, chansync_data_in0_c, chansync_data_in0_d};
assign {chansync_data_out0_de, chansync_data_out0_c, chansync_data_out0_d} = chansync_syncbuffer0_dout;
assign chansync_is_control0 = (~chansync_data_out0_de);
assign chansync_syncbuffer0_re = ((~chansync_is_control0) | chansync_all_control);
assign chansync_syncbuffer1_din = {chansync_data_in1_de, chansync_data_in1_c, chansync_data_in1_d};
assign {chansync_data_out1_de, chansync_data_out1_c, chansync_data_out1_d} = chansync_syncbuffer1_dout;
assign chansync_is_control1 = (~chansync_data_out1_de);
assign chansync_syncbuffer1_re = ((~chansync_is_control1) | chansync_all_control);
assign chansync_syncbuffer2_din = {chansync_data_in2_de, chansync_data_in2_c, chansync_data_in2_d};
assign {chansync_data_out2_de, chansync_data_out2_c, chansync_data_out2_d} = chansync_syncbuffer2_dout;
assign chansync_is_control2 = (~chansync_data_out2_de);
assign chansync_syncbuffer2_re = ((~chansync_is_control2) | chansync_all_control);
assign chansync_all_control = ((chansync_is_control0 & chansync_is_control1) & chansync_is_control2);
assign chansync_some_control = ((chansync_is_control0 | chansync_is_control1) | chansync_is_control2);
assign chansync_syncbuffer0_wrport_adr = chansync_syncbuffer0_produce;
assign chansync_syncbuffer0_wrport_dat_w = chansync_syncbuffer0_din;
assign chansync_syncbuffer0_wrport_we = 1'd1;
assign chansync_syncbuffer0_rdport_adr = chansync_syncbuffer0_consume;
assign chansync_syncbuffer0_dout = chansync_syncbuffer0_rdport_dat_r;
assign chansync_syncbuffer1_wrport_adr = chansync_syncbuffer1_produce;
assign chansync_syncbuffer1_wrport_dat_w = chansync_syncbuffer1_din;
assign chansync_syncbuffer1_wrport_we = 1'd1;
assign chansync_syncbuffer1_rdport_adr = chansync_syncbuffer1_consume;
assign chansync_syncbuffer1_dout = chansync_syncbuffer1_rdport_dat_r;
assign chansync_syncbuffer2_wrport_adr = chansync_syncbuffer2_produce;
assign chansync_syncbuffer2_wrport_dat_w = chansync_syncbuffer2_din;
assign chansync_syncbuffer2_wrport_we = 1'd1;
assign chansync_syncbuffer2_rdport_adr = chansync_syncbuffer2_consume;
assign chansync_syncbuffer2_dout = chansync_syncbuffer2_rdport_dat_r;
assign syncpol_de = syncpol_de_r;
assign syncpol_hsync = syncpol_c_out[0];
assign syncpol_vsync = syncpol_c_out[1];
assign resdetection_pn_de = ((~resdetection_de) & resdetection_de_r);
assign resdetection_p_vsync = (resdetection_vsync & (~resdetection_vsync_r));
assign frame_rgb2ycbcr_sink_valid = frame_valid_i;
assign frame_rgb2ycbcr_sink_payload_r = frame_r;
assign frame_rgb2ycbcr_sink_payload_g = frame_g;
assign frame_rgb2ycbcr_sink_payload_b = frame_b;
assign frame_chroma_downsampler_sink_valid = frame_rgb2ycbcr_source_valid;
assign frame_rgb2ycbcr_source_ready = frame_chroma_downsampler_sink_ready;
assign frame_chroma_downsampler_sink_first = frame_rgb2ycbcr_source_first;
assign frame_chroma_downsampler_sink_last = frame_rgb2ycbcr_source_last;
assign frame_chroma_downsampler_sink_payload_y = frame_rgb2ycbcr_source_payload_y;
assign frame_chroma_downsampler_sink_payload_cb = frame_rgb2ycbcr_source_payload_cb;
assign frame_chroma_downsampler_sink_payload_cr = frame_rgb2ycbcr_source_payload_cr;
assign frame_chroma_downsampler_source_ready = 1'd1;
assign frame_chroma_downsampler_first = (frame_de & (~frame_de_r));
assign frame_new_frame = (frame_next_vsync10 & (~frame_vsync_r));
assign frame_encoded_pixel = {frame_chroma_downsampler_source_payload_cb_cr, frame_chroma_downsampler_source_payload_y};
assign frame_fifo_sink_payload_pixels = frame_cur_word;
assign frame_fifo_sink_valid = frame_cur_word_valid;
assign frame_frame_valid = frame_fifo_source_valid;
assign frame_fifo_source_ready = frame_frame_ready;
assign frame_frame_first = frame_fifo_source_first;
assign frame_frame_last = frame_fifo_source_last;
assign frame_frame_payload_sof = frame_fifo_source_payload_sof;
assign frame_frame_payload_pixels = frame_fifo_source_payload_pixels;
assign frame_busy = 1'd0;
assign frame_pix_overflow_reset = frame_overflow_reset_o;
assign frame_overflow_reset_ack_i = frame_pix_overflow_reset;
assign frame_overflow_w = (frame_sys_overflow & (~frame_overflow_mask));
assign frame_overflow_reset_i = frame_overflow_re;
assign frame_rgb2ycbcr_pipe_ce = (frame_rgb2ycbcr_source_ready | (~frame_rgb2ycbcr_valid_n7));
assign frame_rgb2ycbcr_sink_ready = frame_rgb2ycbcr_pipe_ce;
assign frame_rgb2ycbcr_source_valid = frame_rgb2ycbcr_valid_n7;
assign frame_rgb2ycbcr_busy = ((((((((1'd0 | frame_rgb2ycbcr_valid_n0) | frame_rgb2ycbcr_valid_n1) | frame_rgb2ycbcr_valid_n2) | frame_rgb2ycbcr_valid_n3) | frame_rgb2ycbcr_valid_n4) | frame_rgb2ycbcr_valid_n5) | frame_rgb2ycbcr_valid_n6) | frame_rgb2ycbcr_valid_n7);
assign frame_rgb2ycbcr_source_first = frame_rgb2ycbcr_first_n7;
assign frame_rgb2ycbcr_source_last = frame_rgb2ycbcr_last_n7;
assign frame_rgb2ycbcr_ce = frame_rgb2ycbcr_pipe_ce;
assign frame_rgb2ycbcr_sink_r = frame_rgb2ycbcr_sink_payload_r;
assign frame_rgb2ycbcr_sink_g = frame_rgb2ycbcr_sink_payload_g;
assign frame_rgb2ycbcr_sink_b = frame_rgb2ycbcr_sink_payload_b;
assign frame_rgb2ycbcr_source_payload_y = frame_rgb2ycbcr_source_y;
assign frame_rgb2ycbcr_source_payload_cb = frame_rgb2ycbcr_source_cb;
assign frame_rgb2ycbcr_source_payload_cr = frame_rgb2ycbcr_source_cr;
assign frame_chroma_downsampler_pipe_ce = (frame_chroma_downsampler_source_ready | (~frame_chroma_downsampler_valid_n2));
assign frame_chroma_downsampler_sink_ready = frame_chroma_downsampler_pipe_ce;
assign frame_chroma_downsampler_source_valid = frame_chroma_downsampler_valid_n2;
assign frame_chroma_downsampler_busy = (((1'd0 | frame_chroma_downsampler_valid_n0) | frame_chroma_downsampler_valid_n1) | frame_chroma_downsampler_valid_n2);
assign frame_chroma_downsampler_source_first = frame_chroma_downsampler_first_n2;
assign frame_chroma_downsampler_source_last = frame_chroma_downsampler_last_n2;
assign frame_chroma_downsampler_ce = frame_chroma_downsampler_pipe_ce;
assign frame_chroma_downsampler_sink_y = frame_chroma_downsampler_sink_payload_y;
assign frame_chroma_downsampler_sink_cb = frame_chroma_downsampler_sink_payload_cb;
assign frame_chroma_downsampler_sink_cr = frame_chroma_downsampler_sink_payload_cr;
assign frame_chroma_downsampler_source_payload_y = frame_chroma_downsampler_source_y;
assign frame_chroma_downsampler_source_payload_cb_cr = frame_chroma_downsampler_source_cb_cr;
assign frame_chroma_downsampler_cb_mean = frame_chroma_downsampler_cb_sum[8:1];
assign frame_chroma_downsampler_cr_mean = frame_chroma_downsampler_cr_sum[8:1];
assign frame_fifo_asyncfifo_din = {frame_fifo_fifo_in_last, frame_fifo_fifo_in_first, frame_fifo_fifo_in_payload_pixels, frame_fifo_fifo_in_payload_sof};
assign {frame_fifo_fifo_out_last, frame_fifo_fifo_out_first, frame_fifo_fifo_out_payload_pixels, frame_fifo_fifo_out_payload_sof} = frame_fifo_asyncfifo_dout;
assign frame_fifo_sink_ready = frame_fifo_asyncfifo_writable;
assign frame_fifo_asyncfifo_we = frame_fifo_sink_valid;
assign frame_fifo_fifo_in_first = frame_fifo_sink_first;
assign frame_fifo_fifo_in_last = frame_fifo_sink_last;
assign frame_fifo_fifo_in_payload_sof = frame_fifo_sink_payload_sof;
assign frame_fifo_fifo_in_payload_pixels = frame_fifo_sink_payload_pixels;
assign frame_fifo_source_valid = frame_fifo_asyncfifo_readable;
assign frame_fifo_source_first = frame_fifo_fifo_out_first;
assign frame_fifo_source_last = frame_fifo_fifo_out_last;
assign frame_fifo_source_payload_sof = frame_fifo_fifo_out_payload_sof;
assign frame_fifo_source_payload_pixels = frame_fifo_fifo_out_payload_pixels;
assign frame_fifo_asyncfifo_re = frame_fifo_source_ready;
assign frame_fifo_graycounter0_ce = (frame_fifo_asyncfifo_writable & frame_fifo_asyncfifo_we);
assign frame_fifo_graycounter1_ce = (frame_fifo_asyncfifo_readable & frame_fifo_asyncfifo_re);
assign frame_fifo_asyncfifo_writable = (((frame_fifo_graycounter0_q[9] == frame_fifo_consume_wdomain[9]) | (frame_fifo_graycounter0_q[8] == frame_fifo_consume_wdomain[8])) | (frame_fifo_graycounter0_q[7:0] != frame_fifo_consume_wdomain[7:0]));
assign frame_fifo_asyncfifo_readable = (frame_fifo_graycounter1_q != frame_fifo_produce_rdomain);
assign frame_fifo_wrport_adr = frame_fifo_graycounter0_q_binary[8:0];
assign frame_fifo_wrport_dat_w = frame_fifo_asyncfifo_din;
assign frame_fifo_wrport_we = frame_fifo_graycounter0_ce;
assign frame_fifo_rdport_adr = frame_fifo_graycounter1_q_next_binary[8:0];
assign frame_fifo_asyncfifo_dout = frame_fifo_rdport_dat_r;
always @(*) begin
	frame_fifo_graycounter0_q_next_binary <= 10'd0;
	if (frame_fifo_graycounter0_ce) begin
		frame_fifo_graycounter0_q_next_binary <= (frame_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		frame_fifo_graycounter0_q_next_binary <= frame_fifo_graycounter0_q_binary;
	end
end
assign frame_fifo_graycounter0_q_next = (frame_fifo_graycounter0_q_next_binary ^ frame_fifo_graycounter0_q_next_binary[9:1]);
always @(*) begin
	frame_fifo_graycounter1_q_next_binary <= 10'd0;
	if (frame_fifo_graycounter1_ce) begin
		frame_fifo_graycounter1_q_next_binary <= (frame_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		frame_fifo_graycounter1_q_next_binary <= frame_fifo_graycounter1_q_binary;
	end
end
assign frame_fifo_graycounter1_q_next = (frame_fifo_graycounter1_q_next_binary ^ frame_fifo_graycounter1_q_next_binary[9:1]);
assign frame_overflow_reset_o = (frame_overflow_reset_toggle_o ^ frame_overflow_reset_toggle_o_r);
assign frame_overflow_reset_ack_o = (frame_overflow_reset_ack_toggle_o ^ frame_overflow_reset_ack_toggle_o_r);
assign dma_slot_array_address_reached = dma_current_address;
assign dma_last_word = (dma_mwords_remaining == 1'd1);
assign dma_memory_word = {dma_frame_payload_pixels, dma_frame_payload_pixels, dma_frame_payload_pixels, dma_frame_payload_pixels, dma_frame_payload_pixels, dma_frame_payload_pixels, dma_frame_payload_pixels, dma_frame_payload_pixels};
assign dma_sink_sink_payload_address = dma_current_address;
assign dma_sink_sink_payload_data = dma_memory_word;
assign dma_slot_array_change_slot = ((~dma_slot_array_address_valid) | dma_slot_array_address_done);
assign dma_slot_array_address = comb_rhs_array_muxed36;
assign dma_slot_array_address_valid = comb_rhs_array_muxed37;
assign dma_slot_array_slot0_address_reached = dma_slot_array_address_reached;
assign dma_slot_array_slot1_address_reached = dma_slot_array_address_reached;
assign dma_slot_array_slot0_address_done = (dma_slot_array_address_done & (dma_slot_array_current_slot == 1'd0));
assign dma_slot_array_slot1_address_done = (dma_slot_array_address_done & (dma_slot_array_current_slot == 1'd1));
always @(*) begin
	dma_slot_array_slot0_clear <= 1'd0;
	if ((dma_slot_array_pending_re & dma_slot_array_pending_r[0])) begin
		dma_slot_array_slot0_clear <= 1'd1;
	end
end
always @(*) begin
	dma_slot_array_status_w <= 2'd0;
	dma_slot_array_status_w[0] <= dma_slot_array_slot0_status;
	dma_slot_array_status_w[1] <= dma_slot_array_slot1_status;
end
always @(*) begin
	dma_slot_array_slot1_clear <= 1'd0;
	if ((dma_slot_array_pending_re & dma_slot_array_pending_r[1])) begin
		dma_slot_array_slot1_clear <= 1'd1;
	end
end
always @(*) begin
	dma_slot_array_pending_w <= 2'd0;
	dma_slot_array_pending_w[0] <= dma_slot_array_slot0_pending;
	dma_slot_array_pending_w[1] <= dma_slot_array_slot1_pending;
end
assign dma_slot_array_irq = ((dma_slot_array_pending_w[0] & dma_slot_array_storage[0]) | (dma_slot_array_pending_w[1] & dma_slot_array_storage[1]));
assign dma_slot_array_slot0_status = dma_slot_array_slot0_trigger;
assign dma_slot_array_slot0_pending = dma_slot_array_slot0_trigger;
assign dma_slot_array_slot1_status = dma_slot_array_slot1_trigger;
assign dma_slot_array_slot1_pending = dma_slot_array_slot1_trigger;
assign dma_slot_array_slot0_address = dma_slot_array_slot0_address_storage;
assign dma_slot_array_slot0_address_valid = dma_slot_array_slot0_status_storage[0];
assign dma_slot_array_slot0_status_dat_w = 2'd2;
assign dma_slot_array_slot0_status_we = dma_slot_array_slot0_address_done;
assign dma_slot_array_slot0_address_dat_w = dma_slot_array_slot0_address_reached;
assign dma_slot_array_slot0_address_we = dma_slot_array_slot0_address_done;
assign dma_slot_array_slot0_trigger = dma_slot_array_slot0_status_storage[1];
assign dma_slot_array_slot1_address = dma_slot_array_slot1_address_storage;
assign dma_slot_array_slot1_address_valid = dma_slot_array_slot1_status_storage[0];
assign dma_slot_array_slot1_status_dat_w = 2'd2;
assign dma_slot_array_slot1_status_we = dma_slot_array_slot1_address_done;
assign dma_slot_array_slot1_address_dat_w = dma_slot_array_slot1_address_reached;
assign dma_slot_array_slot1_address_we = dma_slot_array_slot1_address_done;
assign dma_slot_array_slot1_trigger = dma_slot_array_slot1_status_storage[1];
assign litedramcrossbar_cmd_payload_we = 1'd1;
assign litedramcrossbar_cmd_valid = (dma_fifo_sink_ready & dma_sink_sink_valid);
assign litedramcrossbar_cmd_payload_adr = dma_sink_sink_payload_address;
assign dma_sink_sink_ready = (dma_fifo_sink_ready & litedramcrossbar_cmd_ready);
assign dma_fifo_sink_valid = (dma_sink_sink_valid & litedramcrossbar_cmd_ready);
assign dma_fifo_sink_payload_data = dma_sink_sink_payload_data;
assign litedramcrossbar_wdata_valid = dma_fifo_source_valid;
assign dma_fifo_source_ready = litedramcrossbar_wdata_ready;
assign litedramcrossbar_wdata_payload_we = 16'd65535;
assign litedramcrossbar_wdata_payload_data = dma_fifo_source_payload_data;
assign dma_fifo_syncfifo_din = {dma_fifo_fifo_in_last, dma_fifo_fifo_in_first, dma_fifo_fifo_in_payload_data};
assign {dma_fifo_fifo_out_last, dma_fifo_fifo_out_first, dma_fifo_fifo_out_payload_data} = dma_fifo_syncfifo_dout;
assign dma_fifo_sink_ready = dma_fifo_syncfifo_writable;
assign dma_fifo_syncfifo_we = dma_fifo_sink_valid;
assign dma_fifo_fifo_in_first = dma_fifo_sink_first;
assign dma_fifo_fifo_in_last = dma_fifo_sink_last;
assign dma_fifo_fifo_in_payload_data = dma_fifo_sink_payload_data;
assign dma_fifo_source_valid = dma_fifo_syncfifo_readable;
assign dma_fifo_source_first = dma_fifo_fifo_out_first;
assign dma_fifo_source_last = dma_fifo_fifo_out_last;
assign dma_fifo_source_payload_data = dma_fifo_fifo_out_payload_data;
assign dma_fifo_syncfifo_re = dma_fifo_source_ready;
always @(*) begin
	dma_fifo_wrport_adr <= 4'd0;
	if (dma_fifo_replace) begin
		dma_fifo_wrport_adr <= (dma_fifo_produce - 1'd1);
	end else begin
		dma_fifo_wrport_adr <= dma_fifo_produce;
	end
end
assign dma_fifo_wrport_dat_w = dma_fifo_syncfifo_din;
assign dma_fifo_wrport_we = (dma_fifo_syncfifo_we & (dma_fifo_syncfifo_writable | dma_fifo_replace));
assign dma_fifo_do_read = (dma_fifo_syncfifo_readable & dma_fifo_syncfifo_re);
assign dma_fifo_rdport_adr = dma_fifo_consume;
assign dma_fifo_syncfifo_dout = dma_fifo_rdport_dat_r;
assign dma_fifo_syncfifo_writable = (dma_fifo_level != 5'd16);
assign dma_fifo_syncfifo_readable = (dma_fifo_level != 1'd0);
always @(*) begin
	dma_reset_words <= 1'd0;
	dma_count_word <= 1'd0;
	dma_sink_sink_valid <= 1'd0;
	dma_next_state <= 2'd0;
	dma_slot_array_address_done <= 1'd0;
	dma_frame_ready <= 1'd0;
	dma_next_state <= dma_state;
	case (dma_state)
		1'd1: begin
			dma_frame_ready <= dma_sink_sink_ready;
			if (dma_frame_valid) begin
				dma_sink_sink_valid <= 1'd1;
				if (dma_sink_sink_ready) begin
					dma_count_word <= 1'd1;
					if (dma_last_word) begin
						dma_next_state <= 2'd2;
					end
				end
			end
		end
		2'd2: begin
			if ((~litedramcrossbar_wdata_valid)) begin
				dma_slot_array_address_done <= 1'd1;
				dma_next_state <= 1'd0;
			end
		end
		default: begin
			dma_reset_words <= 1'd1;
			dma_frame_ready <= ((~dma_slot_array_address_valid) | (~dma_frame_payload_sof));
			if (((dma_slot_array_address_valid & dma_frame_payload_sof) & dma_frame_valid)) begin
				dma_next_state <= 1'd1;
			end
		end
	endcase
end
assign fmeter_clk = hdmi_in0_freq_clk0;
assign hdmi_in0_freq_period_done = (hdmi_in0_freq_period_counter == 27'd100000000);
assign hdmi_in0_freq_ce = 1'd1;
assign hdmi_in0_freq_sampler_latch = hdmi_in0_freq_period_done;
assign hdmi_in0_freq_sampler_i = hdmi_in0_freq_gray_decoder_o;
assign hdmi_in0_freq_status = hdmi_in0_freq_sampler_o;
always @(*) begin
	hdmi_in0_freq_q_next_binary <= 6'd0;
	if (hdmi_in0_freq_ce) begin
		hdmi_in0_freq_q_next_binary <= (hdmi_in0_freq_q_binary + 1'd1);
	end else begin
		hdmi_in0_freq_q_next_binary <= hdmi_in0_freq_q_binary;
	end
end
assign hdmi_in0_freq_q_next = (hdmi_in0_freq_q_next_binary ^ hdmi_in0_freq_q_next_binary[5:1]);
always @(*) begin
	hdmi_in0_freq_gray_decoder_o_comb <= 6'd0;
	hdmi_in0_freq_gray_decoder_o_comb[5] <= hdmi_in0_freq_gray_decoder_i[5];
	hdmi_in0_freq_gray_decoder_o_comb[4] <= (hdmi_in0_freq_gray_decoder_o_comb[5] ^ hdmi_in0_freq_gray_decoder_i[4]);
	hdmi_in0_freq_gray_decoder_o_comb[3] <= (hdmi_in0_freq_gray_decoder_o_comb[4] ^ hdmi_in0_freq_gray_decoder_i[3]);
	hdmi_in0_freq_gray_decoder_o_comb[2] <= (hdmi_in0_freq_gray_decoder_o_comb[3] ^ hdmi_in0_freq_gray_decoder_i[2]);
	hdmi_in0_freq_gray_decoder_o_comb[1] <= (hdmi_in0_freq_gray_decoder_o_comb[2] ^ hdmi_in0_freq_gray_decoder_i[1]);
	hdmi_in0_freq_gray_decoder_o_comb[0] <= (hdmi_in0_freq_gray_decoder_o_comb[1] ^ hdmi_in0_freq_gray_decoder_i[0]);
end
assign hdmi_in0_freq_sampler_inc = (hdmi_in0_freq_sampler_i - hdmi_in0_freq_sampler_i_d);
assign hdmi_out0_core_source_source_ready = 1'd1;
assign hdmi_out0_resetinserter_reset = (hdmi_out0_core_source_source_param_de & (~hdmi_out0_de_r));
assign hdmi_out0_resetinserter_sink_sink_valid = hdmi_out0_core_source_valid_d;
assign hdmi_out0_resetinserter_sink_sink_payload_y = hdmi_out0_core_source_data_d[7:0];
assign hdmi_out0_resetinserter_sink_sink_payload_cb_cr = hdmi_out0_core_source_data_d[15:8];
assign hdmi_out0_sink_valid = hdmi_out0_resetinserter_source_source_valid;
assign hdmi_out0_resetinserter_source_source_ready = hdmi_out0_sink_ready;
assign hdmi_out0_sink_first = hdmi_out0_resetinserter_source_source_first;
assign hdmi_out0_sink_last = hdmi_out0_resetinserter_source_source_last;
assign hdmi_out0_sink_payload_y = hdmi_out0_resetinserter_source_source_payload_y;
assign hdmi_out0_sink_payload_cb = hdmi_out0_resetinserter_source_source_payload_cb;
assign hdmi_out0_sink_payload_cr = hdmi_out0_resetinserter_source_source_payload_cr;
assign hdmi_out0_driver_sink_sink_valid = hdmi_out0_source_valid;
assign hdmi_out0_source_ready = hdmi_out0_driver_sink_sink_ready;
assign hdmi_out0_driver_sink_sink_first = hdmi_out0_source_first;
assign hdmi_out0_driver_sink_sink_last = hdmi_out0_source_last;
assign hdmi_out0_driver_sink_sink_payload_r = hdmi_out0_source_payload_r;
assign hdmi_out0_driver_sink_sink_payload_g = hdmi_out0_source_payload_g;
assign hdmi_out0_driver_sink_sink_payload_b = hdmi_out0_source_payload_b;
assign hdmi_out0_sink_payload_de = hdmi_out0_core_source_source_param_de;
assign hdmi_out0_sink_payload_vsync = hdmi_out0_core_source_source_param_vsync;
assign hdmi_out0_sink_payload_hsync = hdmi_out0_core_source_source_param_hsync;
assign hdmi_out0_driver_sink_sink_param_de = hdmi_out0_source_payload_de;
assign hdmi_out0_driver_sink_sink_param_vsync = hdmi_out0_source_payload_vsync;
assign hdmi_out0_driver_sink_sink_param_hsync = hdmi_out0_source_payload_hsync;
assign hdmi_out0_core_timinggenerator_sink_valid = hdmi_out0_core_initiator_source_source_valid;
assign hdmi_out0_core_dmareader_sink_valid = hdmi_out0_core_initiator_source_source_valid;
assign hdmi_out0_core_initiator_source_source_ready = hdmi_out0_core_timinggenerator_sink_ready;
assign hdmi_out0_core_source_source_valid = (hdmi_out0_core_timinggenerator_source_valid & ((~hdmi_out0_core_timinggenerator_source_payload_de) | hdmi_out0_core_dmareader_source_valid));
always @(*) begin
	hdmi_out0_core_timinggenerator_source_ready <= 1'd0;
	hdmi_out0_core_dmareader_source_ready <= 1'd0;
	if ((~hdmi_out0_core_initiator_source_source_valid)) begin
		hdmi_out0_core_timinggenerator_source_ready <= 1'd1;
		hdmi_out0_core_dmareader_source_ready <= 1'd1;
	end else begin
		if ((hdmi_out0_core_source_source_valid & hdmi_out0_core_source_source_ready)) begin
			hdmi_out0_core_timinggenerator_source_ready <= 1'd1;
			hdmi_out0_core_dmareader_source_ready <= hdmi_out0_core_timinggenerator_source_payload_de;
		end
	end
end
assign hdmi_out0_core_timinggenerator_sink_payload_hres = hdmi_out0_core_initiator_source_source_payload_hres;
assign hdmi_out0_core_timinggenerator_sink_payload_hsync_start = hdmi_out0_core_initiator_source_source_payload_hsync_start;
assign hdmi_out0_core_timinggenerator_sink_payload_hsync_end = hdmi_out0_core_initiator_source_source_payload_hsync_end;
assign hdmi_out0_core_timinggenerator_sink_payload_hscan = hdmi_out0_core_initiator_source_source_payload_hscan;
assign hdmi_out0_core_timinggenerator_sink_payload_vres = hdmi_out0_core_initiator_source_source_payload_vres;
assign hdmi_out0_core_timinggenerator_sink_payload_vsync_start = hdmi_out0_core_initiator_source_source_payload_vsync_start;
assign hdmi_out0_core_timinggenerator_sink_payload_vsync_end = hdmi_out0_core_initiator_source_source_payload_vsync_end;
assign hdmi_out0_core_timinggenerator_sink_payload_vscan = hdmi_out0_core_initiator_source_source_payload_vscan;
assign hdmi_out0_core_dmareader_sink_payload_base = hdmi_out0_core_initiator_source_source_payload_base;
assign hdmi_out0_core_dmareader_sink_payload_length = hdmi_out0_core_initiator_source_source_payload_length;
assign hdmi_out0_core_source_source_param_de = hdmi_out0_core_timinggenerator_source_payload_de;
assign hdmi_out0_core_source_source_param_hsync = hdmi_out0_core_timinggenerator_source_payload_hsync;
assign hdmi_out0_core_source_source_param_vsync = hdmi_out0_core_timinggenerator_source_payload_vsync;
assign hdmi_out0_core_source_source_payload_data = hdmi_out0_core_dmareader_source_payload_data;
assign hdmi_out0_core_i = hdmi_out0_core_underflow_update_underflow_update_re;
assign hdmi_out0_core_underflow_update = hdmi_out0_core_o;
assign hdmi_out0_core_initiator_cdc_sink_payload_hres = hdmi_out0_core_initiator_csrstorage0_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_hsync_start = hdmi_out0_core_initiator_csrstorage1_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_hsync_end = hdmi_out0_core_initiator_csrstorage2_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_hscan = hdmi_out0_core_initiator_csrstorage3_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_vres = hdmi_out0_core_initiator_csrstorage4_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_vsync_start = hdmi_out0_core_initiator_csrstorage5_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_vsync_end = hdmi_out0_core_initiator_csrstorage6_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_vscan = hdmi_out0_core_initiator_csrstorage7_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_base = hdmi_out0_core_initiator_csrstorage8_storage;
assign hdmi_out0_core_initiator_cdc_sink_payload_length = hdmi_out0_core_initiator_csrstorage9_storage;
assign hdmi_out0_core_initiator_cdc_sink_valid = hdmi_out0_core_initiator_enable_storage;
assign hdmi_out0_core_initiator_source_source_valid = hdmi_out0_core_initiator_cdc_source_valid;
assign hdmi_out0_core_initiator_cdc_source_ready = hdmi_out0_core_initiator_source_source_ready;
assign hdmi_out0_core_initiator_source_source_first = hdmi_out0_core_initiator_cdc_source_first;
assign hdmi_out0_core_initiator_source_source_last = hdmi_out0_core_initiator_cdc_source_last;
assign hdmi_out0_core_initiator_source_source_payload_hres = hdmi_out0_core_initiator_cdc_source_payload_hres;
assign hdmi_out0_core_initiator_source_source_payload_hsync_start = hdmi_out0_core_initiator_cdc_source_payload_hsync_start;
assign hdmi_out0_core_initiator_source_source_payload_hsync_end = hdmi_out0_core_initiator_cdc_source_payload_hsync_end;
assign hdmi_out0_core_initiator_source_source_payload_hscan = hdmi_out0_core_initiator_cdc_source_payload_hscan;
assign hdmi_out0_core_initiator_source_source_payload_vres = hdmi_out0_core_initiator_cdc_source_payload_vres;
assign hdmi_out0_core_initiator_source_source_payload_vsync_start = hdmi_out0_core_initiator_cdc_source_payload_vsync_start;
assign hdmi_out0_core_initiator_source_source_payload_vsync_end = hdmi_out0_core_initiator_cdc_source_payload_vsync_end;
assign hdmi_out0_core_initiator_source_source_payload_vscan = hdmi_out0_core_initiator_cdc_source_payload_vscan;
assign hdmi_out0_core_initiator_source_source_payload_base = hdmi_out0_core_initiator_cdc_source_payload_base;
assign hdmi_out0_core_initiator_source_source_payload_length = hdmi_out0_core_initiator_cdc_source_payload_length;
assign hdmi_out0_core_initiator_cdc_asyncfifo_din = {hdmi_out0_core_initiator_cdc_fifo_in_last, hdmi_out0_core_initiator_cdc_fifo_in_first, hdmi_out0_core_initiator_cdc_fifo_in_payload_length, hdmi_out0_core_initiator_cdc_fifo_in_payload_base, hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan, hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end, hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start, hdmi_out0_core_initiator_cdc_fifo_in_payload_vres, hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan, hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end, hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start, hdmi_out0_core_initiator_cdc_fifo_in_payload_hres};
assign {hdmi_out0_core_initiator_cdc_fifo_out_last, hdmi_out0_core_initiator_cdc_fifo_out_first, hdmi_out0_core_initiator_cdc_fifo_out_payload_length, hdmi_out0_core_initiator_cdc_fifo_out_payload_base, hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan, hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end, hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start, hdmi_out0_core_initiator_cdc_fifo_out_payload_vres, hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan, hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end, hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start, hdmi_out0_core_initiator_cdc_fifo_out_payload_hres} = hdmi_out0_core_initiator_cdc_asyncfifo_dout;
assign hdmi_out0_core_initiator_cdc_sink_ready = hdmi_out0_core_initiator_cdc_asyncfifo_writable;
assign hdmi_out0_core_initiator_cdc_asyncfifo_we = hdmi_out0_core_initiator_cdc_sink_valid;
assign hdmi_out0_core_initiator_cdc_fifo_in_first = hdmi_out0_core_initiator_cdc_sink_first;
assign hdmi_out0_core_initiator_cdc_fifo_in_last = hdmi_out0_core_initiator_cdc_sink_last;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_hres = hdmi_out0_core_initiator_cdc_sink_payload_hres;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start = hdmi_out0_core_initiator_cdc_sink_payload_hsync_start;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end = hdmi_out0_core_initiator_cdc_sink_payload_hsync_end;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan = hdmi_out0_core_initiator_cdc_sink_payload_hscan;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_vres = hdmi_out0_core_initiator_cdc_sink_payload_vres;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start = hdmi_out0_core_initiator_cdc_sink_payload_vsync_start;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end = hdmi_out0_core_initiator_cdc_sink_payload_vsync_end;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan = hdmi_out0_core_initiator_cdc_sink_payload_vscan;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_base = hdmi_out0_core_initiator_cdc_sink_payload_base;
assign hdmi_out0_core_initiator_cdc_fifo_in_payload_length = hdmi_out0_core_initiator_cdc_sink_payload_length;
assign hdmi_out0_core_initiator_cdc_source_valid = hdmi_out0_core_initiator_cdc_asyncfifo_readable;
assign hdmi_out0_core_initiator_cdc_source_first = hdmi_out0_core_initiator_cdc_fifo_out_first;
assign hdmi_out0_core_initiator_cdc_source_last = hdmi_out0_core_initiator_cdc_fifo_out_last;
assign hdmi_out0_core_initiator_cdc_source_payload_hres = hdmi_out0_core_initiator_cdc_fifo_out_payload_hres;
assign hdmi_out0_core_initiator_cdc_source_payload_hsync_start = hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start;
assign hdmi_out0_core_initiator_cdc_source_payload_hsync_end = hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end;
assign hdmi_out0_core_initiator_cdc_source_payload_hscan = hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan;
assign hdmi_out0_core_initiator_cdc_source_payload_vres = hdmi_out0_core_initiator_cdc_fifo_out_payload_vres;
assign hdmi_out0_core_initiator_cdc_source_payload_vsync_start = hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start;
assign hdmi_out0_core_initiator_cdc_source_payload_vsync_end = hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end;
assign hdmi_out0_core_initiator_cdc_source_payload_vscan = hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan;
assign hdmi_out0_core_initiator_cdc_source_payload_base = hdmi_out0_core_initiator_cdc_fifo_out_payload_base;
assign hdmi_out0_core_initiator_cdc_source_payload_length = hdmi_out0_core_initiator_cdc_fifo_out_payload_length;
assign hdmi_out0_core_initiator_cdc_asyncfifo_re = hdmi_out0_core_initiator_cdc_source_ready;
assign hdmi_out0_core_initiator_cdc_graycounter0_ce = (hdmi_out0_core_initiator_cdc_asyncfifo_writable & hdmi_out0_core_initiator_cdc_asyncfifo_we);
assign hdmi_out0_core_initiator_cdc_graycounter1_ce = (hdmi_out0_core_initiator_cdc_asyncfifo_readable & hdmi_out0_core_initiator_cdc_asyncfifo_re);
assign hdmi_out0_core_initiator_cdc_asyncfifo_writable = ((hdmi_out0_core_initiator_cdc_graycounter0_q[1] == hdmi_out0_core_initiator_cdc_consume_wdomain[1]) | (hdmi_out0_core_initiator_cdc_graycounter0_q[0] == hdmi_out0_core_initiator_cdc_consume_wdomain[0]));
assign hdmi_out0_core_initiator_cdc_asyncfifo_readable = (hdmi_out0_core_initiator_cdc_graycounter1_q != hdmi_out0_core_initiator_cdc_produce_rdomain);
assign hdmi_out0_core_initiator_cdc_wrport_adr = hdmi_out0_core_initiator_cdc_graycounter0_q_binary[0];
assign hdmi_out0_core_initiator_cdc_wrport_dat_w = hdmi_out0_core_initiator_cdc_asyncfifo_din;
assign hdmi_out0_core_initiator_cdc_wrport_we = hdmi_out0_core_initiator_cdc_graycounter0_ce;
assign hdmi_out0_core_initiator_cdc_rdport_adr = hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary[0];
assign hdmi_out0_core_initiator_cdc_asyncfifo_dout = hdmi_out0_core_initiator_cdc_rdport_dat_r;
always @(*) begin
	hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= 2'd0;
	if (hdmi_out0_core_initiator_cdc_graycounter0_ce) begin
		hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= (hdmi_out0_core_initiator_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= hdmi_out0_core_initiator_cdc_graycounter0_q_binary;
	end
end
assign hdmi_out0_core_initiator_cdc_graycounter0_q_next = (hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary ^ hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary[1]);
always @(*) begin
	hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= 2'd0;
	if (hdmi_out0_core_initiator_cdc_graycounter1_ce) begin
		hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= (hdmi_out0_core_initiator_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= hdmi_out0_core_initiator_cdc_graycounter1_q_binary;
	end
end
assign hdmi_out0_core_initiator_cdc_graycounter1_q_next = (hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary ^ hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary[1]);
always @(*) begin
	hdmi_out0_core_timinggenerator_active <= 1'd0;
	hdmi_out0_core_timinggenerator_source_payload_de <= 1'd0;
	hdmi_out0_core_timinggenerator_source_valid <= 1'd0;
	if (hdmi_out0_core_timinggenerator_sink_valid) begin
		hdmi_out0_core_timinggenerator_active <= (hdmi_out0_core_timinggenerator_hactive & hdmi_out0_core_timinggenerator_vactive);
		hdmi_out0_core_timinggenerator_source_valid <= 1'd1;
		if (hdmi_out0_core_timinggenerator_active) begin
			hdmi_out0_core_timinggenerator_source_payload_de <= 1'd1;
		end
	end
end
assign hdmi_out0_core_timinggenerator_sink_ready = (hdmi_out0_core_timinggenerator_source_ready & hdmi_out0_core_timinggenerator_source_last);
assign hdmi_out0_core_dmareader_base = hdmi_out0_core_dmareader_sink_payload_base[31:1];
assign hdmi_out0_core_dmareader_length = hdmi_out0_core_dmareader_sink_payload_length[31:1];
assign hdmi_out0_core_dmareader_sink_sink_payload_address = (hdmi_out0_core_dmareader_base + hdmi_out0_core_dmareader_offset);
assign hdmi_out0_core_dmareader_source_valid = hdmi_out0_core_dmareader_source_source_valid;
assign hdmi_out0_core_dmareader_source_source_ready = hdmi_out0_core_dmareader_source_ready;
assign hdmi_out0_core_dmareader_source_first = hdmi_out0_core_dmareader_source_source_first;
assign hdmi_out0_core_dmareader_source_last = hdmi_out0_core_dmareader_source_source_last;
assign hdmi_out0_core_dmareader_source_payload_data = hdmi_out0_core_dmareader_source_source_payload_data;
assign hdmi_out0_dram_port_litedramport1_cmd_payload_we = 1'd0;
assign hdmi_out0_dram_port_litedramport1_cmd_valid = (hdmi_out0_core_dmareader_sink_sink_valid & hdmi_out0_core_dmareader_request_enable);
assign hdmi_out0_dram_port_litedramport1_cmd_payload_adr = hdmi_out0_core_dmareader_sink_sink_payload_address;
assign hdmi_out0_core_dmareader_sink_sink_ready = (hdmi_out0_dram_port_litedramport1_cmd_ready & hdmi_out0_core_dmareader_request_enable);
assign hdmi_out0_core_dmareader_request_issued = (hdmi_out0_dram_port_litedramport1_cmd_valid & hdmi_out0_dram_port_litedramport1_cmd_ready);
assign hdmi_out0_core_dmareader_request_enable = (hdmi_out0_core_dmareader_rsv_level != 13'd4096);
assign hdmi_out0_core_dmareader_fifo_sink_valid = hdmi_out0_dram_port_litedramport1_rdata_valid;
assign hdmi_out0_dram_port_litedramport1_rdata_ready = hdmi_out0_core_dmareader_fifo_sink_ready;
assign hdmi_out0_core_dmareader_fifo_sink_first = hdmi_out0_dram_port_litedramport1_rdata_first;
assign hdmi_out0_core_dmareader_fifo_sink_last = hdmi_out0_dram_port_litedramport1_rdata_last;
assign hdmi_out0_core_dmareader_fifo_sink_payload_data = hdmi_out0_dram_port_litedramport1_rdata_payload_data;
assign hdmi_out0_core_dmareader_source_source_valid = hdmi_out0_core_dmareader_fifo_source_valid;
assign hdmi_out0_core_dmareader_fifo_source_ready = hdmi_out0_core_dmareader_source_source_ready;
assign hdmi_out0_core_dmareader_source_source_first = hdmi_out0_core_dmareader_fifo_source_first;
assign hdmi_out0_core_dmareader_source_source_last = hdmi_out0_core_dmareader_fifo_source_last;
assign hdmi_out0_core_dmareader_source_source_payload_data = hdmi_out0_core_dmareader_fifo_source_payload_data;
assign hdmi_out0_core_dmareader_data_dequeued = (hdmi_out0_core_dmareader_source_source_valid & hdmi_out0_core_dmareader_source_source_ready);
assign hdmi_out0_core_dmareader_fifo_syncfifo_din = {hdmi_out0_core_dmareader_fifo_fifo_in_last, hdmi_out0_core_dmareader_fifo_fifo_in_first, hdmi_out0_core_dmareader_fifo_fifo_in_payload_data};
assign {hdmi_out0_core_dmareader_fifo_fifo_out_last, hdmi_out0_core_dmareader_fifo_fifo_out_first, hdmi_out0_core_dmareader_fifo_fifo_out_payload_data} = hdmi_out0_core_dmareader_fifo_syncfifo_dout;
assign hdmi_out0_core_dmareader_fifo_sink_ready = hdmi_out0_core_dmareader_fifo_syncfifo_writable;
assign hdmi_out0_core_dmareader_fifo_syncfifo_we = hdmi_out0_core_dmareader_fifo_sink_valid;
assign hdmi_out0_core_dmareader_fifo_fifo_in_first = hdmi_out0_core_dmareader_fifo_sink_first;
assign hdmi_out0_core_dmareader_fifo_fifo_in_last = hdmi_out0_core_dmareader_fifo_sink_last;
assign hdmi_out0_core_dmareader_fifo_fifo_in_payload_data = hdmi_out0_core_dmareader_fifo_sink_payload_data;
assign hdmi_out0_core_dmareader_fifo_source_valid = hdmi_out0_core_dmareader_fifo_readable;
assign hdmi_out0_core_dmareader_fifo_source_first = hdmi_out0_core_dmareader_fifo_fifo_out_first;
assign hdmi_out0_core_dmareader_fifo_source_last = hdmi_out0_core_dmareader_fifo_fifo_out_last;
assign hdmi_out0_core_dmareader_fifo_source_payload_data = hdmi_out0_core_dmareader_fifo_fifo_out_payload_data;
assign hdmi_out0_core_dmareader_fifo_re = hdmi_out0_core_dmareader_fifo_source_ready;
assign hdmi_out0_core_dmareader_fifo_syncfifo_re = (hdmi_out0_core_dmareader_fifo_syncfifo_readable & ((~hdmi_out0_core_dmareader_fifo_readable) | hdmi_out0_core_dmareader_fifo_re));
assign hdmi_out0_core_dmareader_fifo_level1 = (hdmi_out0_core_dmareader_fifo_level0 + hdmi_out0_core_dmareader_fifo_readable);
always @(*) begin
	hdmi_out0_core_dmareader_fifo_wrport_adr <= 12'd0;
	if (hdmi_out0_core_dmareader_fifo_replace) begin
		hdmi_out0_core_dmareader_fifo_wrport_adr <= (hdmi_out0_core_dmareader_fifo_produce - 1'd1);
	end else begin
		hdmi_out0_core_dmareader_fifo_wrport_adr <= hdmi_out0_core_dmareader_fifo_produce;
	end
end
assign hdmi_out0_core_dmareader_fifo_wrport_dat_w = hdmi_out0_core_dmareader_fifo_syncfifo_din;
assign hdmi_out0_core_dmareader_fifo_wrport_we = (hdmi_out0_core_dmareader_fifo_syncfifo_we & (hdmi_out0_core_dmareader_fifo_syncfifo_writable | hdmi_out0_core_dmareader_fifo_replace));
assign hdmi_out0_core_dmareader_fifo_do_read = (hdmi_out0_core_dmareader_fifo_syncfifo_readable & hdmi_out0_core_dmareader_fifo_syncfifo_re);
assign hdmi_out0_core_dmareader_fifo_rdport_adr = hdmi_out0_core_dmareader_fifo_consume;
assign hdmi_out0_core_dmareader_fifo_syncfifo_dout = hdmi_out0_core_dmareader_fifo_rdport_dat_r;
assign hdmi_out0_core_dmareader_fifo_rdport_re = hdmi_out0_core_dmareader_fifo_do_read;
assign hdmi_out0_core_dmareader_fifo_syncfifo_writable = (hdmi_out0_core_dmareader_fifo_level0 != 13'd4096);
assign hdmi_out0_core_dmareader_fifo_syncfifo_readable = (hdmi_out0_core_dmareader_fifo_level0 != 1'd0);
always @(*) begin
	hdmi_out0_core_dmareader_sink_sink_valid <= 1'd0;
	hdmi_out0_core_dmareader_offset_videoout_next_value_ce <= 1'd0;
	videoout_next_state <= 1'd0;
	hdmi_out0_core_dmareader_offset_videoout_next_value <= 28'd0;
	hdmi_out0_core_dmareader_sink_ready <= 1'd0;
	hdmi_out0_dram_port_litedramport1_flush <= 1'd0;
	videoout_next_state <= videoout_state;
	case (videoout_state)
		1'd1: begin
			hdmi_out0_core_dmareader_sink_sink_valid <= 1'd1;
			if (hdmi_out0_core_dmareader_sink_sink_ready) begin
				hdmi_out0_core_dmareader_offset_videoout_next_value <= (hdmi_out0_core_dmareader_offset + 1'd1);
				hdmi_out0_core_dmareader_offset_videoout_next_value_ce <= 1'd1;
				if ((hdmi_out0_core_dmareader_offset == (hdmi_out0_core_dmareader_length - 1'd1))) begin
					hdmi_out0_core_dmareader_sink_ready <= 1'd1;
					videoout_next_state <= 1'd0;
				end
			end
		end
		default: begin
			hdmi_out0_core_dmareader_offset_videoout_next_value <= 1'd0;
			hdmi_out0_core_dmareader_offset_videoout_next_value_ce <= 1'd1;
			if (hdmi_out0_core_dmareader_sink_valid) begin
				videoout_next_state <= 1'd1;
			end else begin
				hdmi_out0_dram_port_litedramport1_flush <= 1'd1;
			end
		end
	endcase
end
assign hdmi_out0_core_o = (hdmi_out0_core_toggle_o ^ hdmi_out0_core_toggle_o_r);
assign hdmi_out0_driver_hdmi_phy_sink_valid = hdmi_out0_driver_sink_sink_valid;
assign hdmi_out0_driver_sink_sink_ready = hdmi_out0_driver_hdmi_phy_sink_ready;
assign hdmi_out0_driver_hdmi_phy_sink_first = hdmi_out0_driver_sink_sink_first;
assign hdmi_out0_driver_hdmi_phy_sink_last = hdmi_out0_driver_sink_sink_last;
assign hdmi_out0_driver_hdmi_phy_sink_payload_r = hdmi_out0_driver_sink_sink_payload_r;
assign hdmi_out0_driver_hdmi_phy_sink_payload_g = hdmi_out0_driver_sink_sink_payload_g;
assign hdmi_out0_driver_hdmi_phy_sink_payload_b = hdmi_out0_driver_sink_sink_payload_b;
assign hdmi_out0_driver_hdmi_phy_sink_param_hsync = hdmi_out0_driver_sink_sink_param_hsync;
assign hdmi_out0_driver_hdmi_phy_sink_param_vsync = hdmi_out0_driver_sink_sink_param_vsync;
assign hdmi_out0_driver_hdmi_phy_sink_param_de = hdmi_out0_driver_sink_sink_param_de;
assign hdmi_out0_pix_rst = (~hdmi_out0_driver_s7hdmioutclocking_mmcm_locked);
assign hdmi_out0_driver_s7hdmioutclocking_data0 = hdmi_out0_driver_s7hdmioutclocking;
assign hdmi_out0_driver_s7hdmioutclocking_data1 = hdmi_out0_driver_s7hdmioutclocking_data0;
assign hdmi_out0_driver_hdmi_phy_sink_ready = 1'd1;
assign hdmi_out0_driver_hdmi_phy_es0_d0 = hdmi_out0_driver_hdmi_phy_sink_payload_b;
assign hdmi_out0_driver_hdmi_phy_es1_d0 = hdmi_out0_driver_hdmi_phy_sink_payload_g;
assign hdmi_out0_driver_hdmi_phy_es2_d0 = hdmi_out0_driver_hdmi_phy_sink_payload_r;
assign hdmi_out0_driver_hdmi_phy_es0_c = {hdmi_out0_driver_hdmi_phy_sink_param_vsync, hdmi_out0_driver_hdmi_phy_sink_param_hsync};
assign hdmi_out0_driver_hdmi_phy_es1_c = 1'd0;
assign hdmi_out0_driver_hdmi_phy_es2_c = 1'd0;
assign hdmi_out0_driver_hdmi_phy_es0_de = hdmi_out0_driver_hdmi_phy_sink_param_de;
assign hdmi_out0_driver_hdmi_phy_es1_de = hdmi_out0_driver_hdmi_phy_sink_param_de;
assign hdmi_out0_driver_hdmi_phy_es2_de = hdmi_out0_driver_hdmi_phy_sink_param_de;
assign hdmi_out0_driver_hdmi_phy_es0_data = hdmi_out0_driver_hdmi_phy_es0_out;
assign hdmi_out0_driver_hdmi_phy_es0_q_m8_n = ((hdmi_out0_driver_hdmi_phy_es0_n1d > 3'd4) | ((hdmi_out0_driver_hdmi_phy_es0_n1d == 3'd4) & (~hdmi_out0_driver_hdmi_phy_es0_d1[0])));
assign hdmi_out0_driver_hdmi_phy_es1_data = hdmi_out0_driver_hdmi_phy_es1_out;
assign hdmi_out0_driver_hdmi_phy_es1_q_m8_n = ((hdmi_out0_driver_hdmi_phy_es1_n1d > 3'd4) | ((hdmi_out0_driver_hdmi_phy_es1_n1d == 3'd4) & (~hdmi_out0_driver_hdmi_phy_es1_d1[0])));
assign hdmi_out0_driver_hdmi_phy_es2_data = hdmi_out0_driver_hdmi_phy_es2_out;
assign hdmi_out0_driver_hdmi_phy_es2_q_m8_n = ((hdmi_out0_driver_hdmi_phy_es2_n1d > 3'd4) | ((hdmi_out0_driver_hdmi_phy_es2_n1d == 3'd4) & (~hdmi_out0_driver_hdmi_phy_es2_d1[0])));
always @(*) begin
	hdmi_out0_resetinserter_y_fifo_sink_valid <= 1'd0;
	hdmi_out0_resetinserter_cb_fifo_sink_valid <= 1'd0;
	hdmi_out0_resetinserter_cr_fifo_sink_valid <= 1'd0;
	hdmi_out0_resetinserter_y_fifo_sink_payload_data <= 8'd0;
	hdmi_out0_resetinserter_cb_fifo_sink_payload_data <= 8'd0;
	hdmi_out0_resetinserter_cr_fifo_sink_payload_data <= 8'd0;
	hdmi_out0_resetinserter_sink_sink_ready <= 1'd0;
	if ((~hdmi_out0_resetinserter_parity_in)) begin
		hdmi_out0_resetinserter_y_fifo_sink_valid <= (hdmi_out0_resetinserter_sink_sink_valid & hdmi_out0_resetinserter_sink_sink_ready);
		hdmi_out0_resetinserter_y_fifo_sink_payload_data <= hdmi_out0_resetinserter_sink_sink_payload_y;
		hdmi_out0_resetinserter_cb_fifo_sink_valid <= (hdmi_out0_resetinserter_sink_sink_valid & hdmi_out0_resetinserter_sink_sink_ready);
		hdmi_out0_resetinserter_cb_fifo_sink_payload_data <= hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
		hdmi_out0_resetinserter_sink_sink_ready <= (hdmi_out0_resetinserter_y_fifo_sink_ready & hdmi_out0_resetinserter_cb_fifo_sink_ready);
	end else begin
		hdmi_out0_resetinserter_y_fifo_sink_valid <= (hdmi_out0_resetinserter_sink_sink_valid & hdmi_out0_resetinserter_sink_sink_ready);
		hdmi_out0_resetinserter_y_fifo_sink_payload_data <= hdmi_out0_resetinserter_sink_sink_payload_y;
		hdmi_out0_resetinserter_cr_fifo_sink_valid <= (hdmi_out0_resetinserter_sink_sink_valid & hdmi_out0_resetinserter_sink_sink_ready);
		hdmi_out0_resetinserter_cr_fifo_sink_payload_data <= hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
		hdmi_out0_resetinserter_sink_sink_ready <= (hdmi_out0_resetinserter_y_fifo_sink_ready & hdmi_out0_resetinserter_cr_fifo_sink_ready);
	end
end
assign hdmi_out0_resetinserter_source_source_valid = ((hdmi_out0_resetinserter_y_fifo_source_valid & hdmi_out0_resetinserter_cb_fifo_source_valid) & hdmi_out0_resetinserter_cr_fifo_source_valid);
assign hdmi_out0_resetinserter_source_source_payload_y = hdmi_out0_resetinserter_y_fifo_source_payload_data;
assign hdmi_out0_resetinserter_source_source_payload_cb = hdmi_out0_resetinserter_cb_fifo_source_payload_data;
assign hdmi_out0_resetinserter_source_source_payload_cr = hdmi_out0_resetinserter_cr_fifo_source_payload_data;
assign hdmi_out0_resetinserter_y_fifo_source_ready = (hdmi_out0_resetinserter_source_source_valid & hdmi_out0_resetinserter_source_source_ready);
assign hdmi_out0_resetinserter_cb_fifo_source_ready = ((hdmi_out0_resetinserter_source_source_valid & hdmi_out0_resetinserter_source_source_ready) & hdmi_out0_resetinserter_parity_out);
assign hdmi_out0_resetinserter_cr_fifo_source_ready = ((hdmi_out0_resetinserter_source_source_valid & hdmi_out0_resetinserter_source_source_ready) & hdmi_out0_resetinserter_parity_out);
assign hdmi_out0_resetinserter_y_fifo_syncfifo_din = {hdmi_out0_resetinserter_y_fifo_fifo_in_last, hdmi_out0_resetinserter_y_fifo_fifo_in_first, hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data};
assign {hdmi_out0_resetinserter_y_fifo_fifo_out_last, hdmi_out0_resetinserter_y_fifo_fifo_out_first, hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data} = hdmi_out0_resetinserter_y_fifo_syncfifo_dout;
assign hdmi_out0_resetinserter_y_fifo_sink_ready = hdmi_out0_resetinserter_y_fifo_syncfifo_writable;
assign hdmi_out0_resetinserter_y_fifo_syncfifo_we = hdmi_out0_resetinserter_y_fifo_sink_valid;
assign hdmi_out0_resetinserter_y_fifo_fifo_in_first = hdmi_out0_resetinserter_y_fifo_sink_first;
assign hdmi_out0_resetinserter_y_fifo_fifo_in_last = hdmi_out0_resetinserter_y_fifo_sink_last;
assign hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data = hdmi_out0_resetinserter_y_fifo_sink_payload_data;
assign hdmi_out0_resetinserter_y_fifo_source_valid = hdmi_out0_resetinserter_y_fifo_syncfifo_readable;
assign hdmi_out0_resetinserter_y_fifo_source_first = hdmi_out0_resetinserter_y_fifo_fifo_out_first;
assign hdmi_out0_resetinserter_y_fifo_source_last = hdmi_out0_resetinserter_y_fifo_fifo_out_last;
assign hdmi_out0_resetinserter_y_fifo_source_payload_data = hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data;
assign hdmi_out0_resetinserter_y_fifo_syncfifo_re = hdmi_out0_resetinserter_y_fifo_source_ready;
always @(*) begin
	hdmi_out0_resetinserter_y_fifo_wrport_adr <= 2'd0;
	if (hdmi_out0_resetinserter_y_fifo_replace) begin
		hdmi_out0_resetinserter_y_fifo_wrport_adr <= (hdmi_out0_resetinserter_y_fifo_produce - 1'd1);
	end else begin
		hdmi_out0_resetinserter_y_fifo_wrport_adr <= hdmi_out0_resetinserter_y_fifo_produce;
	end
end
assign hdmi_out0_resetinserter_y_fifo_wrport_dat_w = hdmi_out0_resetinserter_y_fifo_syncfifo_din;
assign hdmi_out0_resetinserter_y_fifo_wrport_we = (hdmi_out0_resetinserter_y_fifo_syncfifo_we & (hdmi_out0_resetinserter_y_fifo_syncfifo_writable | hdmi_out0_resetinserter_y_fifo_replace));
assign hdmi_out0_resetinserter_y_fifo_do_read = (hdmi_out0_resetinserter_y_fifo_syncfifo_readable & hdmi_out0_resetinserter_y_fifo_syncfifo_re);
assign hdmi_out0_resetinserter_y_fifo_rdport_adr = hdmi_out0_resetinserter_y_fifo_consume;
assign hdmi_out0_resetinserter_y_fifo_syncfifo_dout = hdmi_out0_resetinserter_y_fifo_rdport_dat_r;
assign hdmi_out0_resetinserter_y_fifo_syncfifo_writable = (hdmi_out0_resetinserter_y_fifo_level != 3'd4);
assign hdmi_out0_resetinserter_y_fifo_syncfifo_readable = (hdmi_out0_resetinserter_y_fifo_level != 1'd0);
assign hdmi_out0_resetinserter_cb_fifo_syncfifo_din = {hdmi_out0_resetinserter_cb_fifo_fifo_in_last, hdmi_out0_resetinserter_cb_fifo_fifo_in_first, hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data};
assign {hdmi_out0_resetinserter_cb_fifo_fifo_out_last, hdmi_out0_resetinserter_cb_fifo_fifo_out_first, hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data} = hdmi_out0_resetinserter_cb_fifo_syncfifo_dout;
assign hdmi_out0_resetinserter_cb_fifo_sink_ready = hdmi_out0_resetinserter_cb_fifo_syncfifo_writable;
assign hdmi_out0_resetinserter_cb_fifo_syncfifo_we = hdmi_out0_resetinserter_cb_fifo_sink_valid;
assign hdmi_out0_resetinserter_cb_fifo_fifo_in_first = hdmi_out0_resetinserter_cb_fifo_sink_first;
assign hdmi_out0_resetinserter_cb_fifo_fifo_in_last = hdmi_out0_resetinserter_cb_fifo_sink_last;
assign hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data = hdmi_out0_resetinserter_cb_fifo_sink_payload_data;
assign hdmi_out0_resetinserter_cb_fifo_source_valid = hdmi_out0_resetinserter_cb_fifo_syncfifo_readable;
assign hdmi_out0_resetinserter_cb_fifo_source_first = hdmi_out0_resetinserter_cb_fifo_fifo_out_first;
assign hdmi_out0_resetinserter_cb_fifo_source_last = hdmi_out0_resetinserter_cb_fifo_fifo_out_last;
assign hdmi_out0_resetinserter_cb_fifo_source_payload_data = hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data;
assign hdmi_out0_resetinserter_cb_fifo_syncfifo_re = hdmi_out0_resetinserter_cb_fifo_source_ready;
always @(*) begin
	hdmi_out0_resetinserter_cb_fifo_wrport_adr <= 2'd0;
	if (hdmi_out0_resetinserter_cb_fifo_replace) begin
		hdmi_out0_resetinserter_cb_fifo_wrport_adr <= (hdmi_out0_resetinserter_cb_fifo_produce - 1'd1);
	end else begin
		hdmi_out0_resetinserter_cb_fifo_wrport_adr <= hdmi_out0_resetinserter_cb_fifo_produce;
	end
end
assign hdmi_out0_resetinserter_cb_fifo_wrport_dat_w = hdmi_out0_resetinserter_cb_fifo_syncfifo_din;
assign hdmi_out0_resetinserter_cb_fifo_wrport_we = (hdmi_out0_resetinserter_cb_fifo_syncfifo_we & (hdmi_out0_resetinserter_cb_fifo_syncfifo_writable | hdmi_out0_resetinserter_cb_fifo_replace));
assign hdmi_out0_resetinserter_cb_fifo_do_read = (hdmi_out0_resetinserter_cb_fifo_syncfifo_readable & hdmi_out0_resetinserter_cb_fifo_syncfifo_re);
assign hdmi_out0_resetinserter_cb_fifo_rdport_adr = hdmi_out0_resetinserter_cb_fifo_consume;
assign hdmi_out0_resetinserter_cb_fifo_syncfifo_dout = hdmi_out0_resetinserter_cb_fifo_rdport_dat_r;
assign hdmi_out0_resetinserter_cb_fifo_syncfifo_writable = (hdmi_out0_resetinserter_cb_fifo_level != 3'd4);
assign hdmi_out0_resetinserter_cb_fifo_syncfifo_readable = (hdmi_out0_resetinserter_cb_fifo_level != 1'd0);
assign hdmi_out0_resetinserter_cr_fifo_syncfifo_din = {hdmi_out0_resetinserter_cr_fifo_fifo_in_last, hdmi_out0_resetinserter_cr_fifo_fifo_in_first, hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data};
assign {hdmi_out0_resetinserter_cr_fifo_fifo_out_last, hdmi_out0_resetinserter_cr_fifo_fifo_out_first, hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data} = hdmi_out0_resetinserter_cr_fifo_syncfifo_dout;
assign hdmi_out0_resetinserter_cr_fifo_sink_ready = hdmi_out0_resetinserter_cr_fifo_syncfifo_writable;
assign hdmi_out0_resetinserter_cr_fifo_syncfifo_we = hdmi_out0_resetinserter_cr_fifo_sink_valid;
assign hdmi_out0_resetinserter_cr_fifo_fifo_in_first = hdmi_out0_resetinserter_cr_fifo_sink_first;
assign hdmi_out0_resetinserter_cr_fifo_fifo_in_last = hdmi_out0_resetinserter_cr_fifo_sink_last;
assign hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data = hdmi_out0_resetinserter_cr_fifo_sink_payload_data;
assign hdmi_out0_resetinserter_cr_fifo_source_valid = hdmi_out0_resetinserter_cr_fifo_syncfifo_readable;
assign hdmi_out0_resetinserter_cr_fifo_source_first = hdmi_out0_resetinserter_cr_fifo_fifo_out_first;
assign hdmi_out0_resetinserter_cr_fifo_source_last = hdmi_out0_resetinserter_cr_fifo_fifo_out_last;
assign hdmi_out0_resetinserter_cr_fifo_source_payload_data = hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data;
assign hdmi_out0_resetinserter_cr_fifo_syncfifo_re = hdmi_out0_resetinserter_cr_fifo_source_ready;
always @(*) begin
	hdmi_out0_resetinserter_cr_fifo_wrport_adr <= 2'd0;
	if (hdmi_out0_resetinserter_cr_fifo_replace) begin
		hdmi_out0_resetinserter_cr_fifo_wrport_adr <= (hdmi_out0_resetinserter_cr_fifo_produce - 1'd1);
	end else begin
		hdmi_out0_resetinserter_cr_fifo_wrport_adr <= hdmi_out0_resetinserter_cr_fifo_produce;
	end
end
assign hdmi_out0_resetinserter_cr_fifo_wrport_dat_w = hdmi_out0_resetinserter_cr_fifo_syncfifo_din;
assign hdmi_out0_resetinserter_cr_fifo_wrport_we = (hdmi_out0_resetinserter_cr_fifo_syncfifo_we & (hdmi_out0_resetinserter_cr_fifo_syncfifo_writable | hdmi_out0_resetinserter_cr_fifo_replace));
assign hdmi_out0_resetinserter_cr_fifo_do_read = (hdmi_out0_resetinserter_cr_fifo_syncfifo_readable & hdmi_out0_resetinserter_cr_fifo_syncfifo_re);
assign hdmi_out0_resetinserter_cr_fifo_rdport_adr = hdmi_out0_resetinserter_cr_fifo_consume;
assign hdmi_out0_resetinserter_cr_fifo_syncfifo_dout = hdmi_out0_resetinserter_cr_fifo_rdport_dat_r;
assign hdmi_out0_resetinserter_cr_fifo_syncfifo_writable = (hdmi_out0_resetinserter_cr_fifo_level != 3'd4);
assign hdmi_out0_resetinserter_cr_fifo_syncfifo_readable = (hdmi_out0_resetinserter_cr_fifo_level != 1'd0);
assign hdmi_out0_pipe_ce = (hdmi_out0_source_ready | (~hdmi_out0_valid_n3));
assign hdmi_out0_sink_ready = hdmi_out0_pipe_ce;
assign hdmi_out0_source_valid = hdmi_out0_valid_n3;
assign hdmi_out0_busy = ((((1'd0 | hdmi_out0_valid_n0) | hdmi_out0_valid_n1) | hdmi_out0_valid_n2) | hdmi_out0_valid_n3);
assign hdmi_out0_source_first = hdmi_out0_first_n3;
assign hdmi_out0_source_last = hdmi_out0_last_n3;
assign hdmi_out0_ce = hdmi_out0_pipe_ce;
assign hdmi_out0_sink_y = hdmi_out0_sink_payload_y;
assign hdmi_out0_sink_cb = hdmi_out0_sink_payload_cb;
assign hdmi_out0_sink_cr = hdmi_out0_sink_payload_cr;
assign hdmi_out0_source_payload_r = hdmi_out0_source_r;
assign hdmi_out0_source_payload_g = hdmi_out0_source_g;
assign hdmi_out0_source_payload_b = hdmi_out0_source_b;
assign hdmi_out0_source_payload_hsync = hdmi_out0_next_s5;
assign hdmi_out0_source_payload_vsync = hdmi_out0_next_s11;
assign hdmi_out0_source_payload_de = hdmi_out0_next_s17;
assign videosoc_interface0_wb_sdram_adr = comb_rhs_array_muxed38;
assign videosoc_interface0_wb_sdram_dat_w = comb_rhs_array_muxed39;
assign videosoc_interface0_wb_sdram_sel = comb_rhs_array_muxed40;
assign videosoc_interface0_wb_sdram_cyc = comb_rhs_array_muxed41;
assign videosoc_interface0_wb_sdram_stb = comb_rhs_array_muxed42;
assign videosoc_interface0_wb_sdram_we = comb_rhs_array_muxed43;
assign videosoc_interface0_wb_sdram_cti = comb_rhs_array_muxed44;
assign videosoc_interface0_wb_sdram_bte = comb_rhs_array_muxed45;
assign videosoc_interface1_wb_sdram_dat_r = videosoc_interface0_wb_sdram_dat_r;
assign videosoc_interface1_wb_sdram_ack = (videosoc_interface0_wb_sdram_ack & (wb_sdram_con_grant == 1'd0));
assign videosoc_interface1_wb_sdram_err = (videosoc_interface0_wb_sdram_err & (wb_sdram_con_grant == 1'd0));
assign wb_sdram_con_request = {videosoc_interface1_wb_sdram_cyc};
assign wb_sdram_con_grant = 1'd0;
assign videosoc_shared_adr = comb_rhs_array_muxed46;
assign videosoc_shared_dat_w = comb_rhs_array_muxed47;
assign videosoc_shared_sel = comb_rhs_array_muxed48;
assign videosoc_shared_cyc = comb_rhs_array_muxed49;
assign videosoc_shared_stb = comb_rhs_array_muxed50;
assign videosoc_shared_we = comb_rhs_array_muxed51;
assign videosoc_shared_cti = comb_rhs_array_muxed52;
assign videosoc_shared_bte = comb_rhs_array_muxed53;
assign videosoc_videosoc_ibus_dat_r = videosoc_shared_dat_r;
assign videosoc_videosoc_dbus_dat_r = videosoc_shared_dat_r;
assign videosoc_bridge_wishbone_dat_r = videosoc_shared_dat_r;
assign videosoc_videosoc_ibus_ack = (videosoc_shared_ack & (videosoc_grant == 1'd0));
assign videosoc_videosoc_dbus_ack = (videosoc_shared_ack & (videosoc_grant == 1'd1));
assign videosoc_bridge_wishbone_ack = (videosoc_shared_ack & (videosoc_grant == 2'd2));
assign videosoc_videosoc_ibus_err = (videosoc_shared_err & (videosoc_grant == 1'd0));
assign videosoc_videosoc_dbus_err = (videosoc_shared_err & (videosoc_grant == 1'd1));
assign videosoc_bridge_wishbone_err = (videosoc_shared_err & (videosoc_grant == 2'd2));
assign videosoc_request = {videosoc_bridge_wishbone_cyc, videosoc_videosoc_dbus_cyc, videosoc_videosoc_ibus_cyc};
always @(*) begin
	videosoc_slave_sel <= 6'd0;
	videosoc_slave_sel[0] <= (videosoc_shared_adr[28:26] == 1'd0);
	videosoc_slave_sel[1] <= (videosoc_shared_adr[28:26] == 1'd1);
	videosoc_slave_sel[2] <= (videosoc_shared_adr[28:26] == 3'd6);
	videosoc_slave_sel[3] <= (videosoc_shared_adr[28:26] == 3'd4);
	videosoc_slave_sel[4] <= (videosoc_shared_adr[28:26] == 2'd2);
	videosoc_slave_sel[5] <= (videosoc_shared_adr[28:26] == 2'd3);
end
assign videosoc_videosoc_rom_bus_adr = videosoc_shared_adr;
assign videosoc_videosoc_rom_bus_dat_w = videosoc_shared_dat_w;
assign videosoc_videosoc_rom_bus_sel = videosoc_shared_sel;
assign videosoc_videosoc_rom_bus_stb = videosoc_shared_stb;
assign videosoc_videosoc_rom_bus_we = videosoc_shared_we;
assign videosoc_videosoc_rom_bus_cti = videosoc_shared_cti;
assign videosoc_videosoc_rom_bus_bte = videosoc_shared_bte;
assign videosoc_videosoc_sram_bus_adr = videosoc_shared_adr;
assign videosoc_videosoc_sram_bus_dat_w = videosoc_shared_dat_w;
assign videosoc_videosoc_sram_bus_sel = videosoc_shared_sel;
assign videosoc_videosoc_sram_bus_stb = videosoc_shared_stb;
assign videosoc_videosoc_sram_bus_we = videosoc_shared_we;
assign videosoc_videosoc_sram_bus_cti = videosoc_shared_cti;
assign videosoc_videosoc_sram_bus_bte = videosoc_shared_bte;
assign videosoc_videosoc_bus_wishbone_adr = videosoc_shared_adr;
assign videosoc_videosoc_bus_wishbone_dat_w = videosoc_shared_dat_w;
assign videosoc_videosoc_bus_wishbone_sel = videosoc_shared_sel;
assign videosoc_videosoc_bus_wishbone_stb = videosoc_shared_stb;
assign videosoc_videosoc_bus_wishbone_we = videosoc_shared_we;
assign videosoc_videosoc_bus_wishbone_cti = videosoc_shared_cti;
assign videosoc_videosoc_bus_wishbone_bte = videosoc_shared_bte;
assign videosoc_interface1_wb_sdram_adr = videosoc_shared_adr;
assign videosoc_interface1_wb_sdram_dat_w = videosoc_shared_dat_w;
assign videosoc_interface1_wb_sdram_sel = videosoc_shared_sel;
assign videosoc_interface1_wb_sdram_stb = videosoc_shared_stb;
assign videosoc_interface1_wb_sdram_we = videosoc_shared_we;
assign videosoc_interface1_wb_sdram_cti = videosoc_shared_cti;
assign videosoc_interface1_wb_sdram_bte = videosoc_shared_bte;
assign videosoc_bus_adr = videosoc_shared_adr;
assign videosoc_bus_dat_w = videosoc_shared_dat_w;
assign videosoc_bus_sel = videosoc_shared_sel;
assign videosoc_bus_stb = videosoc_shared_stb;
assign videosoc_bus_we = videosoc_shared_we;
assign videosoc_bus_cti = videosoc_shared_cti;
assign videosoc_bus_bte = videosoc_shared_bte;
assign ethmac_bus_adr = videosoc_shared_adr;
assign ethmac_bus_dat_w = videosoc_shared_dat_w;
assign ethmac_bus_sel = videosoc_shared_sel;
assign ethmac_bus_stb = videosoc_shared_stb;
assign ethmac_bus_we = videosoc_shared_we;
assign ethmac_bus_cti = videosoc_shared_cti;
assign ethmac_bus_bte = videosoc_shared_bte;
assign videosoc_videosoc_rom_bus_cyc = (videosoc_shared_cyc & videosoc_slave_sel[0]);
assign videosoc_videosoc_sram_bus_cyc = (videosoc_shared_cyc & videosoc_slave_sel[1]);
assign videosoc_videosoc_bus_wishbone_cyc = (videosoc_shared_cyc & videosoc_slave_sel[2]);
assign videosoc_interface1_wb_sdram_cyc = (videosoc_shared_cyc & videosoc_slave_sel[3]);
assign videosoc_bus_cyc = (videosoc_shared_cyc & videosoc_slave_sel[4]);
assign ethmac_bus_cyc = (videosoc_shared_cyc & videosoc_slave_sel[5]);
assign videosoc_shared_ack = (((((videosoc_videosoc_rom_bus_ack | videosoc_videosoc_sram_bus_ack) | videosoc_videosoc_bus_wishbone_ack) | videosoc_interface1_wb_sdram_ack) | videosoc_bus_ack) | ethmac_bus_ack);
assign videosoc_shared_err = (((((videosoc_videosoc_rom_bus_err | videosoc_videosoc_sram_bus_err) | videosoc_videosoc_bus_wishbone_err) | videosoc_interface1_wb_sdram_err) | videosoc_bus_err) | ethmac_bus_err);
assign videosoc_shared_dat_r = (((((({32{videosoc_slave_sel_r[0]}} & videosoc_videosoc_rom_bus_dat_r) | ({32{videosoc_slave_sel_r[1]}} & videosoc_videosoc_sram_bus_dat_r)) | ({32{videosoc_slave_sel_r[2]}} & videosoc_videosoc_bus_wishbone_dat_r)) | ({32{videosoc_slave_sel_r[3]}} & videosoc_interface1_wb_sdram_dat_r)) | ({32{videosoc_slave_sel_r[4]}} & videosoc_bus_dat_r)) | ({32{videosoc_slave_sel_r[5]}} & ethmac_bus_dat_r));
assign videosoc_csrbank0_sel = (videosoc_interface0_bank_bus_adr[13:9] == 4'd11);
assign videosoc_csrbank0_dly_sel0_r = videosoc_interface0_bank_bus_dat_w[1:0];
assign videosoc_csrbank0_dly_sel0_re = ((videosoc_csrbank0_sel & videosoc_interface0_bank_bus_we) & (videosoc_interface0_bank_bus_adr[1:0] == 1'd0));
assign videosoc_ddrphy_rdly_dq_rst_r = videosoc_interface0_bank_bus_dat_w[0];
assign videosoc_ddrphy_rdly_dq_rst_re = ((videosoc_csrbank0_sel & videosoc_interface0_bank_bus_we) & (videosoc_interface0_bank_bus_adr[1:0] == 1'd1));
assign videosoc_ddrphy_rdly_dq_inc_r = videosoc_interface0_bank_bus_dat_w[0];
assign videosoc_ddrphy_rdly_dq_inc_re = ((videosoc_csrbank0_sel & videosoc_interface0_bank_bus_we) & (videosoc_interface0_bank_bus_adr[1:0] == 2'd2));
assign videosoc_ddrphy_rdly_dq_bitslip_r = videosoc_interface0_bank_bus_dat_w[0];
assign videosoc_ddrphy_rdly_dq_bitslip_re = ((videosoc_csrbank0_sel & videosoc_interface0_bank_bus_we) & (videosoc_interface0_bank_bus_adr[1:0] == 2'd3));
assign videosoc_ddrphy_storage = videosoc_ddrphy_storage_full[1:0];
assign videosoc_csrbank0_dly_sel0_w = videosoc_ddrphy_storage_full[1:0];
assign videosoc_csrbank1_sel = (videosoc_interface1_bank_bus_adr[13:9] == 4'd15);
assign videosoc_csrbank1_sram_writer_slot_r = videosoc_interface1_bank_bus_dat_w[0];
assign videosoc_csrbank1_sram_writer_slot_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 1'd0));
assign videosoc_csrbank1_sram_writer_length3_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_length3_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 1'd1));
assign videosoc_csrbank1_sram_writer_length2_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_length2_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 2'd2));
assign videosoc_csrbank1_sram_writer_length1_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_length1_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 2'd3));
assign videosoc_csrbank1_sram_writer_length0_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_length0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 3'd4));
assign videosoc_csrbank1_sram_writer_errors3_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_errors3_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 3'd5));
assign videosoc_csrbank1_sram_writer_errors2_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_errors2_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 3'd6));
assign videosoc_csrbank1_sram_writer_errors1_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_errors1_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 3'd7));
assign videosoc_csrbank1_sram_writer_errors0_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_writer_errors0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd8));
assign ethmac_writer_status_r = videosoc_interface1_bank_bus_dat_w[0];
assign ethmac_writer_status_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd9));
assign ethmac_writer_pending_r = videosoc_interface1_bank_bus_dat_w[0];
assign ethmac_writer_pending_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd10));
assign videosoc_csrbank1_sram_writer_ev_enable0_r = videosoc_interface1_bank_bus_dat_w[0];
assign videosoc_csrbank1_sram_writer_ev_enable0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd11));
assign ethmac_reader_start_r = videosoc_interface1_bank_bus_dat_w[0];
assign ethmac_reader_start_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd12));
assign videosoc_csrbank1_sram_reader_ready_r = videosoc_interface1_bank_bus_dat_w[0];
assign videosoc_csrbank1_sram_reader_ready_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd13));
assign videosoc_csrbank1_sram_reader_level_r = videosoc_interface1_bank_bus_dat_w[1:0];
assign videosoc_csrbank1_sram_reader_level_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd14));
assign videosoc_csrbank1_sram_reader_slot0_r = videosoc_interface1_bank_bus_dat_w[0];
assign videosoc_csrbank1_sram_reader_slot0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 4'd15));
assign videosoc_csrbank1_sram_reader_length1_r = videosoc_interface1_bank_bus_dat_w[2:0];
assign videosoc_csrbank1_sram_reader_length1_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd16));
assign videosoc_csrbank1_sram_reader_length0_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_sram_reader_length0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd17));
assign ethmac_reader_eventmanager_status_r = videosoc_interface1_bank_bus_dat_w[0];
assign ethmac_reader_eventmanager_status_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd18));
assign ethmac_reader_eventmanager_pending_r = videosoc_interface1_bank_bus_dat_w[0];
assign ethmac_reader_eventmanager_pending_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd19));
assign videosoc_csrbank1_sram_reader_ev_enable0_r = videosoc_interface1_bank_bus_dat_w[0];
assign videosoc_csrbank1_sram_reader_ev_enable0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd20));
assign videosoc_csrbank1_preamble_crc_r = videosoc_interface1_bank_bus_dat_w[0];
assign videosoc_csrbank1_preamble_crc_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd21));
assign videosoc_csrbank1_preamble_errors3_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_preamble_errors3_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd22));
assign videosoc_csrbank1_preamble_errors2_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_preamble_errors2_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd23));
assign videosoc_csrbank1_preamble_errors1_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_preamble_errors1_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd24));
assign videosoc_csrbank1_preamble_errors0_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_preamble_errors0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd25));
assign videosoc_csrbank1_crc_errors3_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_crc_errors3_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd26));
assign videosoc_csrbank1_crc_errors2_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_crc_errors2_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd27));
assign videosoc_csrbank1_crc_errors1_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_crc_errors1_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd28));
assign videosoc_csrbank1_crc_errors0_r = videosoc_interface1_bank_bus_dat_w[7:0];
assign videosoc_csrbank1_crc_errors0_re = ((videosoc_csrbank1_sel & videosoc_interface1_bank_bus_we) & (videosoc_interface1_bank_bus_adr[4:0] == 5'd29));
assign videosoc_csrbank1_sram_writer_slot_w = ethmac_writer_slot_status;
assign videosoc_csrbank1_sram_writer_length3_w = ethmac_writer_length_status[31:24];
assign videosoc_csrbank1_sram_writer_length2_w = ethmac_writer_length_status[23:16];
assign videosoc_csrbank1_sram_writer_length1_w = ethmac_writer_length_status[15:8];
assign videosoc_csrbank1_sram_writer_length0_w = ethmac_writer_length_status[7:0];
assign videosoc_csrbank1_sram_writer_errors3_w = ethmac_writer_errors_status[31:24];
assign videosoc_csrbank1_sram_writer_errors2_w = ethmac_writer_errors_status[23:16];
assign videosoc_csrbank1_sram_writer_errors1_w = ethmac_writer_errors_status[15:8];
assign videosoc_csrbank1_sram_writer_errors0_w = ethmac_writer_errors_status[7:0];
assign ethmac_writer_storage = ethmac_writer_storage_full;
assign videosoc_csrbank1_sram_writer_ev_enable0_w = ethmac_writer_storage_full;
assign videosoc_csrbank1_sram_reader_ready_w = ethmac_reader_ready_status;
assign videosoc_csrbank1_sram_reader_level_w = ethmac_reader_level_status[1:0];
assign ethmac_reader_slot_storage = ethmac_reader_slot_storage_full;
assign videosoc_csrbank1_sram_reader_slot0_w = ethmac_reader_slot_storage_full;
assign ethmac_reader_length_storage = ethmac_reader_length_storage_full[10:0];
assign videosoc_csrbank1_sram_reader_length1_w = ethmac_reader_length_storage_full[10:8];
assign videosoc_csrbank1_sram_reader_length0_w = ethmac_reader_length_storage_full[7:0];
assign ethmac_reader_eventmanager_storage = ethmac_reader_eventmanager_storage_full;
assign videosoc_csrbank1_sram_reader_ev_enable0_w = ethmac_reader_eventmanager_storage_full;
assign videosoc_csrbank1_preamble_crc_w = ethmac_preamble_crc_status;
assign videosoc_csrbank1_preamble_errors3_w = ethmac_preamble_errors_status[31:24];
assign videosoc_csrbank1_preamble_errors2_w = ethmac_preamble_errors_status[23:16];
assign videosoc_csrbank1_preamble_errors1_w = ethmac_preamble_errors_status[15:8];
assign videosoc_csrbank1_preamble_errors0_w = ethmac_preamble_errors_status[7:0];
assign videosoc_csrbank1_crc_errors3_w = ethmac_crc_errors_status[31:24];
assign videosoc_csrbank1_crc_errors2_w = ethmac_crc_errors_status[23:16];
assign videosoc_csrbank1_crc_errors1_w = ethmac_crc_errors_status[15:8];
assign videosoc_csrbank1_crc_errors0_w = ethmac_crc_errors_status[7:0];
assign videosoc_csrbank2_sel = (videosoc_interface2_bank_bus_adr[13:9] == 4'd14);
assign videosoc_csrbank2_crg_reset0_r = videosoc_interface2_bank_bus_dat_w[0];
assign videosoc_csrbank2_crg_reset0_re = ((videosoc_csrbank2_sel & videosoc_interface2_bank_bus_we) & (videosoc_interface2_bank_bus_adr[1:0] == 1'd0));
assign videosoc_csrbank2_mdio_w0_r = videosoc_interface2_bank_bus_dat_w[2:0];
assign videosoc_csrbank2_mdio_w0_re = ((videosoc_csrbank2_sel & videosoc_interface2_bank_bus_we) & (videosoc_interface2_bank_bus_adr[1:0] == 1'd1));
assign videosoc_csrbank2_mdio_r_r = videosoc_interface2_bank_bus_dat_w[0];
assign videosoc_csrbank2_mdio_r_re = ((videosoc_csrbank2_sel & videosoc_interface2_bank_bus_we) & (videosoc_interface2_bank_bus_adr[1:0] == 2'd2));
assign ethphy_reset_storage = ethphy_reset_storage_full;
assign videosoc_csrbank2_crg_reset0_w = ethphy_reset_storage_full;
assign ethphy_storage = ethphy_storage_full[2:0];
assign videosoc_csrbank2_mdio_w0_w = ethphy_storage_full[2:0];
assign videosoc_csrbank2_mdio_r_w = ethphy_status;
assign videosoc_sram0_sel = (videosoc_interface0_sram_bus_adr[13:9] == 5'd19);
always @(*) begin
	videosoc_interface0_sram_bus_dat_r <= 8'd0;
	if (videosoc_sram0_sel_r) begin
		videosoc_interface0_sram_bus_dat_r <= videosoc_sram0_dat_r;
	end
end
assign videosoc_sram0_we = (videosoc_sram0_sel & videosoc_interface0_sram_bus_we);
assign videosoc_sram0_dat_w = videosoc_interface0_sram_bus_dat_w;
assign videosoc_sram0_adr = videosoc_interface0_sram_bus_adr[6:0];
assign videosoc_csrbank3_sel = (videosoc_interface3_bank_bus_adr[13:9] == 5'd17);
assign videosoc_csrbank3_edid_hpd_notif_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_edid_hpd_notif_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 1'd0));
assign videosoc_csrbank3_edid_hpd_en0_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_edid_hpd_en0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 1'd1));
assign videosoc_csrbank3_clocking_mmcm_reset0_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_clocking_mmcm_reset0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 2'd2));
assign videosoc_csrbank3_clocking_locked_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_clocking_locked_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 2'd3));
assign mmcm_read_r = videosoc_interface3_bank_bus_dat_w[0];
assign mmcm_read_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 3'd4));
assign mmcm_write_r = videosoc_interface3_bank_bus_dat_w[0];
assign mmcm_write_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 3'd5));
assign videosoc_csrbank3_clocking_mmcm_drdy_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_clocking_mmcm_drdy_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 3'd6));
assign videosoc_csrbank3_clocking_mmcm_adr0_r = videosoc_interface3_bank_bus_dat_w[6:0];
assign videosoc_csrbank3_clocking_mmcm_adr0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 3'd7));
assign videosoc_csrbank3_clocking_mmcm_dat_w1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_clocking_mmcm_dat_w1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd8));
assign videosoc_csrbank3_clocking_mmcm_dat_w0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_clocking_mmcm_dat_w0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd9));
assign videosoc_csrbank3_clocking_mmcm_dat_r1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_clocking_mmcm_dat_r1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd10));
assign videosoc_csrbank3_clocking_mmcm_dat_r0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_clocking_mmcm_dat_r0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd11));
assign s7datacapture0_dly_ctl_r = videosoc_interface3_bank_bus_dat_w[4:0];
assign s7datacapture0_dly_ctl_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd12));
assign videosoc_csrbank3_data0_cap_phase_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign videosoc_csrbank3_data0_cap_phase_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd13));
assign s7datacapture0_phase_reset_r = videosoc_interface3_bank_bus_dat_w[0];
assign s7datacapture0_phase_reset_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd14));
assign videosoc_csrbank3_data0_charsync_char_synced_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_data0_charsync_char_synced_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 4'd15));
assign videosoc_csrbank3_data0_charsync_ctl_pos_r = videosoc_interface3_bank_bus_dat_w[3:0];
assign videosoc_csrbank3_data0_charsync_ctl_pos_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd16));
assign wer0_update_r = videosoc_interface3_bank_bus_dat_w[0];
assign wer0_update_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd17));
assign videosoc_csrbank3_data0_wer_value2_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data0_wer_value2_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd18));
assign videosoc_csrbank3_data0_wer_value1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data0_wer_value1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd19));
assign videosoc_csrbank3_data0_wer_value0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data0_wer_value0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd20));
assign s7datacapture1_dly_ctl_r = videosoc_interface3_bank_bus_dat_w[4:0];
assign s7datacapture1_dly_ctl_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd21));
assign videosoc_csrbank3_data1_cap_phase_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign videosoc_csrbank3_data1_cap_phase_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd22));
assign s7datacapture1_phase_reset_r = videosoc_interface3_bank_bus_dat_w[0];
assign s7datacapture1_phase_reset_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd23));
assign videosoc_csrbank3_data1_charsync_char_synced_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_data1_charsync_char_synced_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd24));
assign videosoc_csrbank3_data1_charsync_ctl_pos_r = videosoc_interface3_bank_bus_dat_w[3:0];
assign videosoc_csrbank3_data1_charsync_ctl_pos_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd25));
assign wer1_update_r = videosoc_interface3_bank_bus_dat_w[0];
assign wer1_update_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd26));
assign videosoc_csrbank3_data1_wer_value2_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data1_wer_value2_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd27));
assign videosoc_csrbank3_data1_wer_value1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data1_wer_value1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd28));
assign videosoc_csrbank3_data1_wer_value0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data1_wer_value0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd29));
assign s7datacapture2_dly_ctl_r = videosoc_interface3_bank_bus_dat_w[4:0];
assign s7datacapture2_dly_ctl_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd30));
assign videosoc_csrbank3_data2_cap_phase_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign videosoc_csrbank3_data2_cap_phase_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 5'd31));
assign s7datacapture2_phase_reset_r = videosoc_interface3_bank_bus_dat_w[0];
assign s7datacapture2_phase_reset_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd32));
assign videosoc_csrbank3_data2_charsync_char_synced_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_data2_charsync_char_synced_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd33));
assign videosoc_csrbank3_data2_charsync_ctl_pos_r = videosoc_interface3_bank_bus_dat_w[3:0];
assign videosoc_csrbank3_data2_charsync_ctl_pos_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd34));
assign wer2_update_r = videosoc_interface3_bank_bus_dat_w[0];
assign wer2_update_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd35));
assign videosoc_csrbank3_data2_wer_value2_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data2_wer_value2_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd36));
assign videosoc_csrbank3_data2_wer_value1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data2_wer_value1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd37));
assign videosoc_csrbank3_data2_wer_value0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_data2_wer_value0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd38));
assign videosoc_csrbank3_chansync_channels_synced_r = videosoc_interface3_bank_bus_dat_w[0];
assign videosoc_csrbank3_chansync_channels_synced_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd39));
assign videosoc_csrbank3_resdetection_hres1_r = videosoc_interface3_bank_bus_dat_w[2:0];
assign videosoc_csrbank3_resdetection_hres1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd40));
assign videosoc_csrbank3_resdetection_hres0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_resdetection_hres0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd41));
assign videosoc_csrbank3_resdetection_vres1_r = videosoc_interface3_bank_bus_dat_w[2:0];
assign videosoc_csrbank3_resdetection_vres1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd42));
assign videosoc_csrbank3_resdetection_vres0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_resdetection_vres0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd43));
assign frame_overflow_r = videosoc_interface3_bank_bus_dat_w[0];
assign frame_overflow_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd44));
assign videosoc_csrbank3_dma_frame_size3_r = videosoc_interface3_bank_bus_dat_w[4:0];
assign videosoc_csrbank3_dma_frame_size3_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd45));
assign videosoc_csrbank3_dma_frame_size2_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_frame_size2_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd46));
assign videosoc_csrbank3_dma_frame_size1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_frame_size1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd47));
assign videosoc_csrbank3_dma_frame_size0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_frame_size0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd48));
assign videosoc_csrbank3_dma_slot0_status0_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign videosoc_csrbank3_dma_slot0_status0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd49));
assign videosoc_csrbank3_dma_slot0_address3_r = videosoc_interface3_bank_bus_dat_w[4:0];
assign videosoc_csrbank3_dma_slot0_address3_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd50));
assign videosoc_csrbank3_dma_slot0_address2_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_slot0_address2_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd51));
assign videosoc_csrbank3_dma_slot0_address1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_slot0_address1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd52));
assign videosoc_csrbank3_dma_slot0_address0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_slot0_address0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd53));
assign videosoc_csrbank3_dma_slot1_status0_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign videosoc_csrbank3_dma_slot1_status0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd54));
assign videosoc_csrbank3_dma_slot1_address3_r = videosoc_interface3_bank_bus_dat_w[4:0];
assign videosoc_csrbank3_dma_slot1_address3_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd55));
assign videosoc_csrbank3_dma_slot1_address2_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_slot1_address2_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd56));
assign videosoc_csrbank3_dma_slot1_address1_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_slot1_address1_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd57));
assign videosoc_csrbank3_dma_slot1_address0_r = videosoc_interface3_bank_bus_dat_w[7:0];
assign videosoc_csrbank3_dma_slot1_address0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd58));
assign dma_slot_array_status_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign dma_slot_array_status_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd59));
assign dma_slot_array_pending_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign dma_slot_array_pending_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd60));
assign videosoc_csrbank3_dma_ev_enable0_r = videosoc_interface3_bank_bus_dat_w[1:0];
assign videosoc_csrbank3_dma_ev_enable0_re = ((videosoc_csrbank3_sel & videosoc_interface3_bank_bus_we) & (videosoc_interface3_bank_bus_adr[5:0] == 6'd61));
assign videosoc_csrbank3_edid_hpd_notif_w = edid_status;
assign edid_storage = edid_storage_full;
assign videosoc_csrbank3_edid_hpd_en0_w = edid_storage_full;
assign mmcm_reset_storage = mmcm_reset_storage_full;
assign videosoc_csrbank3_clocking_mmcm_reset0_w = mmcm_reset_storage_full;
assign videosoc_csrbank3_clocking_locked_w = locked_status;
assign videosoc_csrbank3_clocking_mmcm_drdy_w = mmcm_drdy_status;
assign mmcm_adr_storage = mmcm_adr_storage_full[6:0];
assign videosoc_csrbank3_clocking_mmcm_adr0_w = mmcm_adr_storage_full[6:0];
assign mmcm_dat_w_storage = mmcm_dat_w_storage_full[15:0];
assign videosoc_csrbank3_clocking_mmcm_dat_w1_w = mmcm_dat_w_storage_full[15:8];
assign videosoc_csrbank3_clocking_mmcm_dat_w0_w = mmcm_dat_w_storage_full[7:0];
assign videosoc_csrbank3_clocking_mmcm_dat_r1_w = mmcm_dat_r_status[15:8];
assign videosoc_csrbank3_clocking_mmcm_dat_r0_w = mmcm_dat_r_status[7:0];
assign videosoc_csrbank3_data0_cap_phase_w = s7datacapture0_status[1:0];
assign videosoc_csrbank3_data0_charsync_char_synced_w = charsync0_char_synced_status;
assign videosoc_csrbank3_data0_charsync_ctl_pos_w = charsync0_ctl_pos_status[3:0];
assign videosoc_csrbank3_data0_wer_value2_w = wer0_status[23:16];
assign videosoc_csrbank3_data0_wer_value1_w = wer0_status[15:8];
assign videosoc_csrbank3_data0_wer_value0_w = wer0_status[7:0];
assign videosoc_csrbank3_data1_cap_phase_w = s7datacapture1_status[1:0];
assign videosoc_csrbank3_data1_charsync_char_synced_w = charsync1_char_synced_status;
assign videosoc_csrbank3_data1_charsync_ctl_pos_w = charsync1_ctl_pos_status[3:0];
assign videosoc_csrbank3_data1_wer_value2_w = wer1_status[23:16];
assign videosoc_csrbank3_data1_wer_value1_w = wer1_status[15:8];
assign videosoc_csrbank3_data1_wer_value0_w = wer1_status[7:0];
assign videosoc_csrbank3_data2_cap_phase_w = s7datacapture2_status[1:0];
assign videosoc_csrbank3_data2_charsync_char_synced_w = charsync2_char_synced_status;
assign videosoc_csrbank3_data2_charsync_ctl_pos_w = charsync2_ctl_pos_status[3:0];
assign videosoc_csrbank3_data2_wer_value2_w = wer2_status[23:16];
assign videosoc_csrbank3_data2_wer_value1_w = wer2_status[15:8];
assign videosoc_csrbank3_data2_wer_value0_w = wer2_status[7:0];
assign videosoc_csrbank3_chansync_channels_synced_w = chansync_status;
assign videosoc_csrbank3_resdetection_hres1_w = resdetection_hres_status[10:8];
assign videosoc_csrbank3_resdetection_hres0_w = resdetection_hres_status[7:0];
assign videosoc_csrbank3_resdetection_vres1_w = resdetection_vres_status[10:8];
assign videosoc_csrbank3_resdetection_vres0_w = resdetection_vres_status[7:0];
assign dma_frame_size_storage = dma_frame_size_storage_full[28:4];
assign videosoc_csrbank3_dma_frame_size3_w = dma_frame_size_storage_full[28:24];
assign videosoc_csrbank3_dma_frame_size2_w = dma_frame_size_storage_full[23:16];
assign videosoc_csrbank3_dma_frame_size1_w = dma_frame_size_storage_full[15:8];
assign videosoc_csrbank3_dma_frame_size0_w = {dma_frame_size_storage_full[7:4], {4{1'd0}}};
assign dma_slot_array_slot0_status_storage = dma_slot_array_slot0_status_storage_full[1:0];
assign videosoc_csrbank3_dma_slot0_status0_w = dma_slot_array_slot0_status_storage_full[1:0];
assign dma_slot_array_slot0_address_storage = dma_slot_array_slot0_address_storage_full[28:4];
assign videosoc_csrbank3_dma_slot0_address3_w = dma_slot_array_slot0_address_storage_full[28:24];
assign videosoc_csrbank3_dma_slot0_address2_w = dma_slot_array_slot0_address_storage_full[23:16];
assign videosoc_csrbank3_dma_slot0_address1_w = dma_slot_array_slot0_address_storage_full[15:8];
assign videosoc_csrbank3_dma_slot0_address0_w = {dma_slot_array_slot0_address_storage_full[7:4], {4{1'd0}}};
assign dma_slot_array_slot1_status_storage = dma_slot_array_slot1_status_storage_full[1:0];
assign videosoc_csrbank3_dma_slot1_status0_w = dma_slot_array_slot1_status_storage_full[1:0];
assign dma_slot_array_slot1_address_storage = dma_slot_array_slot1_address_storage_full[28:4];
assign videosoc_csrbank3_dma_slot1_address3_w = dma_slot_array_slot1_address_storage_full[28:24];
assign videosoc_csrbank3_dma_slot1_address2_w = dma_slot_array_slot1_address_storage_full[23:16];
assign videosoc_csrbank3_dma_slot1_address1_w = dma_slot_array_slot1_address_storage_full[15:8];
assign videosoc_csrbank3_dma_slot1_address0_w = {dma_slot_array_slot1_address_storage_full[7:4], {4{1'd0}}};
assign dma_slot_array_storage = dma_slot_array_storage_full[1:0];
assign videosoc_csrbank3_dma_ev_enable0_w = dma_slot_array_storage_full[1:0];
assign videosoc_csrbank4_sel = (videosoc_interface4_bank_bus_adr[13:9] == 5'd18);
assign videosoc_csrbank4_value3_r = videosoc_interface4_bank_bus_dat_w[7:0];
assign videosoc_csrbank4_value3_re = ((videosoc_csrbank4_sel & videosoc_interface4_bank_bus_we) & (videosoc_interface4_bank_bus_adr[1:0] == 1'd0));
assign videosoc_csrbank4_value2_r = videosoc_interface4_bank_bus_dat_w[7:0];
assign videosoc_csrbank4_value2_re = ((videosoc_csrbank4_sel & videosoc_interface4_bank_bus_we) & (videosoc_interface4_bank_bus_adr[1:0] == 1'd1));
assign videosoc_csrbank4_value1_r = videosoc_interface4_bank_bus_dat_w[7:0];
assign videosoc_csrbank4_value1_re = ((videosoc_csrbank4_sel & videosoc_interface4_bank_bus_we) & (videosoc_interface4_bank_bus_adr[1:0] == 2'd2));
assign videosoc_csrbank4_value0_r = videosoc_interface4_bank_bus_dat_w[7:0];
assign videosoc_csrbank4_value0_re = ((videosoc_csrbank4_sel & videosoc_interface4_bank_bus_we) & (videosoc_interface4_bank_bus_adr[1:0] == 2'd3));
assign videosoc_csrbank4_value3_w = hdmi_in0_freq_status[31:24];
assign videosoc_csrbank4_value2_w = hdmi_in0_freq_status[23:16];
assign videosoc_csrbank4_value1_w = hdmi_in0_freq_status[15:8];
assign videosoc_csrbank4_value0_w = hdmi_in0_freq_status[7:0];
assign videosoc_csrbank5_sel = (videosoc_interface5_bank_bus_adr[13:9] == 5'd16);
assign videosoc_csrbank5_core_underflow_enable0_r = videosoc_interface5_bank_bus_dat_w[0];
assign videosoc_csrbank5_core_underflow_enable0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 1'd0));
assign hdmi_out0_core_underflow_update_underflow_update_r = videosoc_interface5_bank_bus_dat_w[0];
assign hdmi_out0_core_underflow_update_underflow_update_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 1'd1));
assign videosoc_csrbank5_core_underflow_counter3_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_underflow_counter3_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 2'd2));
assign videosoc_csrbank5_core_underflow_counter2_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_underflow_counter2_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 2'd3));
assign videosoc_csrbank5_core_underflow_counter1_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_underflow_counter1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 3'd4));
assign videosoc_csrbank5_core_underflow_counter0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_underflow_counter0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 3'd5));
assign videosoc_csrbank5_core_initiator_enable0_r = videosoc_interface5_bank_bus_dat_w[0];
assign videosoc_csrbank5_core_initiator_enable0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 3'd6));
assign videosoc_csrbank5_core_initiator_hres1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_hres1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 3'd7));
assign videosoc_csrbank5_core_initiator_hres0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_hres0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd8));
assign videosoc_csrbank5_core_initiator_hsync_start1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_hsync_start1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd9));
assign videosoc_csrbank5_core_initiator_hsync_start0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_hsync_start0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd10));
assign videosoc_csrbank5_core_initiator_hsync_end1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_hsync_end1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd11));
assign videosoc_csrbank5_core_initiator_hsync_end0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_hsync_end0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd12));
assign videosoc_csrbank5_core_initiator_hscan1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_hscan1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd13));
assign videosoc_csrbank5_core_initiator_hscan0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_hscan0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd14));
assign videosoc_csrbank5_core_initiator_vres1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_vres1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 4'd15));
assign videosoc_csrbank5_core_initiator_vres0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_vres0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd16));
assign videosoc_csrbank5_core_initiator_vsync_start1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_vsync_start1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd17));
assign videosoc_csrbank5_core_initiator_vsync_start0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_vsync_start0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd18));
assign videosoc_csrbank5_core_initiator_vsync_end1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_vsync_end1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd19));
assign videosoc_csrbank5_core_initiator_vsync_end0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_vsync_end0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd20));
assign videosoc_csrbank5_core_initiator_vscan1_r = videosoc_interface5_bank_bus_dat_w[3:0];
assign videosoc_csrbank5_core_initiator_vscan1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd21));
assign videosoc_csrbank5_core_initiator_vscan0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_vscan0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd22));
assign videosoc_csrbank5_core_initiator_base3_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_base3_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd23));
assign videosoc_csrbank5_core_initiator_base2_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_base2_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd24));
assign videosoc_csrbank5_core_initiator_base1_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_base1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd25));
assign videosoc_csrbank5_core_initiator_base0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_base0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd26));
assign videosoc_csrbank5_core_initiator_length3_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_length3_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd27));
assign videosoc_csrbank5_core_initiator_length2_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_length2_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd28));
assign videosoc_csrbank5_core_initiator_length1_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_length1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd29));
assign videosoc_csrbank5_core_initiator_length0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_core_initiator_length0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd30));
assign videosoc_csrbank5_driver_clocking_mmcm_reset0_r = videosoc_interface5_bank_bus_dat_w[0];
assign videosoc_csrbank5_driver_clocking_mmcm_reset0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 5'd31));
assign hdmi_out0_driver_s7hdmioutclocking_mmcm_read_r = videosoc_interface5_bank_bus_dat_w[0];
assign hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd32));
assign hdmi_out0_driver_s7hdmioutclocking_mmcm_write_r = videosoc_interface5_bank_bus_dat_w[0];
assign hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd33));
assign videosoc_csrbank5_driver_clocking_mmcm_drdy_r = videosoc_interface5_bank_bus_dat_w[0];
assign videosoc_csrbank5_driver_clocking_mmcm_drdy_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd34));
assign videosoc_csrbank5_driver_clocking_mmcm_adr0_r = videosoc_interface5_bank_bus_dat_w[6:0];
assign videosoc_csrbank5_driver_clocking_mmcm_adr0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd35));
assign videosoc_csrbank5_driver_clocking_mmcm_dat_w1_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_w1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd36));
assign videosoc_csrbank5_driver_clocking_mmcm_dat_w0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd37));
assign videosoc_csrbank5_driver_clocking_mmcm_dat_r1_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_r1_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd38));
assign videosoc_csrbank5_driver_clocking_mmcm_dat_r0_r = videosoc_interface5_bank_bus_dat_w[7:0];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_r0_re = ((videosoc_csrbank5_sel & videosoc_interface5_bank_bus_we) & (videosoc_interface5_bank_bus_adr[5:0] == 6'd39));
assign hdmi_out0_core_underflow_enable_storage = hdmi_out0_core_underflow_enable_storage_full;
assign videosoc_csrbank5_core_underflow_enable0_w = hdmi_out0_core_underflow_enable_storage_full;
assign videosoc_csrbank5_core_underflow_counter3_w = hdmi_out0_core_underflow_counter_status[31:24];
assign videosoc_csrbank5_core_underflow_counter2_w = hdmi_out0_core_underflow_counter_status[23:16];
assign videosoc_csrbank5_core_underflow_counter1_w = hdmi_out0_core_underflow_counter_status[15:8];
assign videosoc_csrbank5_core_underflow_counter0_w = hdmi_out0_core_underflow_counter_status[7:0];
assign hdmi_out0_core_initiator_enable_storage = hdmi_out0_core_initiator_enable_storage_full;
assign videosoc_csrbank5_core_initiator_enable0_w = hdmi_out0_core_initiator_enable_storage_full;
assign hdmi_out0_core_initiator_csrstorage0_storage = hdmi_out0_core_initiator_csrstorage0_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_hres1_w = hdmi_out0_core_initiator_csrstorage0_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_hres0_w = hdmi_out0_core_initiator_csrstorage0_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage1_storage = hdmi_out0_core_initiator_csrstorage1_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_hsync_start1_w = hdmi_out0_core_initiator_csrstorage1_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_hsync_start0_w = hdmi_out0_core_initiator_csrstorage1_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage2_storage = hdmi_out0_core_initiator_csrstorage2_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_hsync_end1_w = hdmi_out0_core_initiator_csrstorage2_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_hsync_end0_w = hdmi_out0_core_initiator_csrstorage2_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage3_storage = hdmi_out0_core_initiator_csrstorage3_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_hscan1_w = hdmi_out0_core_initiator_csrstorage3_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_hscan0_w = hdmi_out0_core_initiator_csrstorage3_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage4_storage = hdmi_out0_core_initiator_csrstorage4_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_vres1_w = hdmi_out0_core_initiator_csrstorage4_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_vres0_w = hdmi_out0_core_initiator_csrstorage4_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage5_storage = hdmi_out0_core_initiator_csrstorage5_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_vsync_start1_w = hdmi_out0_core_initiator_csrstorage5_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_vsync_start0_w = hdmi_out0_core_initiator_csrstorage5_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage6_storage = hdmi_out0_core_initiator_csrstorage6_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_vsync_end1_w = hdmi_out0_core_initiator_csrstorage6_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_vsync_end0_w = hdmi_out0_core_initiator_csrstorage6_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage7_storage = hdmi_out0_core_initiator_csrstorage7_storage_full[11:0];
assign videosoc_csrbank5_core_initiator_vscan1_w = hdmi_out0_core_initiator_csrstorage7_storage_full[11:8];
assign videosoc_csrbank5_core_initiator_vscan0_w = hdmi_out0_core_initiator_csrstorage7_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage8_storage = hdmi_out0_core_initiator_csrstorage8_storage_full[31:0];
assign videosoc_csrbank5_core_initiator_base3_w = hdmi_out0_core_initiator_csrstorage8_storage_full[31:24];
assign videosoc_csrbank5_core_initiator_base2_w = hdmi_out0_core_initiator_csrstorage8_storage_full[23:16];
assign videosoc_csrbank5_core_initiator_base1_w = hdmi_out0_core_initiator_csrstorage8_storage_full[15:8];
assign videosoc_csrbank5_core_initiator_base0_w = hdmi_out0_core_initiator_csrstorage8_storage_full[7:0];
assign hdmi_out0_core_initiator_csrstorage9_storage = hdmi_out0_core_initiator_csrstorage9_storage_full[31:0];
assign videosoc_csrbank5_core_initiator_length3_w = hdmi_out0_core_initiator_csrstorage9_storage_full[31:24];
assign videosoc_csrbank5_core_initiator_length2_w = hdmi_out0_core_initiator_csrstorage9_storage_full[23:16];
assign videosoc_csrbank5_core_initiator_length1_w = hdmi_out0_core_initiator_csrstorage9_storage_full[15:8];
assign videosoc_csrbank5_core_initiator_length0_w = hdmi_out0_core_initiator_csrstorage9_storage_full[7:0];
assign hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage = hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full;
assign videosoc_csrbank5_driver_clocking_mmcm_reset0_w = hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full;
assign videosoc_csrbank5_driver_clocking_mmcm_drdy_w = hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status;
assign hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage = hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full[6:0];
assign videosoc_csrbank5_driver_clocking_mmcm_adr0_w = hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full[6:0];
assign hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage = hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[15:0];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_w1_w = hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[15:8];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_w0_w = hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[7:0];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_r1_w = hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status[15:8];
assign videosoc_csrbank5_driver_clocking_mmcm_dat_r0_w = hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status[7:0];
assign videosoc_sram1_sel = (videosoc_interface1_sram_bus_adr[13:9] == 2'd3);
always @(*) begin
	videosoc_interface1_sram_bus_dat_r <= 8'd0;
	if (videosoc_sram1_sel_r) begin
		videosoc_interface1_sram_bus_dat_r <= videosoc_sram1_dat_r;
	end
end
assign videosoc_sram1_adr = videosoc_interface1_sram_bus_adr[3:0];
assign videosoc_csrbank6_sel = (videosoc_interface6_bank_bus_adr[13:9] == 4'd12);
assign videosoc_csrbank6_dna_id7_r = videosoc_interface6_bank_bus_dat_w[0];
assign videosoc_csrbank6_dna_id7_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 1'd0));
assign videosoc_csrbank6_dna_id6_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_dna_id6_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 1'd1));
assign videosoc_csrbank6_dna_id5_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_dna_id5_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 2'd2));
assign videosoc_csrbank6_dna_id4_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_dna_id4_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 2'd3));
assign videosoc_csrbank6_dna_id3_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_dna_id3_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 3'd4));
assign videosoc_csrbank6_dna_id2_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_dna_id2_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 3'd5));
assign videosoc_csrbank6_dna_id1_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_dna_id1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 3'd6));
assign videosoc_csrbank6_dna_id0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_dna_id0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 3'd7));
assign videosoc_csrbank6_git_commit19_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit19_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd8));
assign videosoc_csrbank6_git_commit18_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit18_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd9));
assign videosoc_csrbank6_git_commit17_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit17_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd10));
assign videosoc_csrbank6_git_commit16_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit16_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd11));
assign videosoc_csrbank6_git_commit15_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit15_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd12));
assign videosoc_csrbank6_git_commit14_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit14_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd13));
assign videosoc_csrbank6_git_commit13_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit13_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd14));
assign videosoc_csrbank6_git_commit12_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit12_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 4'd15));
assign videosoc_csrbank6_git_commit11_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit11_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd16));
assign videosoc_csrbank6_git_commit10_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit10_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd17));
assign videosoc_csrbank6_git_commit9_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit9_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd18));
assign videosoc_csrbank6_git_commit8_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit8_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd19));
assign videosoc_csrbank6_git_commit7_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit7_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd20));
assign videosoc_csrbank6_git_commit6_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit6_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd21));
assign videosoc_csrbank6_git_commit5_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit5_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd22));
assign videosoc_csrbank6_git_commit4_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit4_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd23));
assign videosoc_csrbank6_git_commit3_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit3_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd24));
assign videosoc_csrbank6_git_commit2_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit2_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd25));
assign videosoc_csrbank6_git_commit1_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd26));
assign videosoc_csrbank6_git_commit0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_git_commit0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd27));
assign videosoc_csrbank6_platform_platform7_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform7_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd28));
assign videosoc_csrbank6_platform_platform6_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform6_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd29));
assign videosoc_csrbank6_platform_platform5_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform5_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd30));
assign videosoc_csrbank6_platform_platform4_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform4_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 5'd31));
assign videosoc_csrbank6_platform_platform3_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform3_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd32));
assign videosoc_csrbank6_platform_platform2_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform2_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd33));
assign videosoc_csrbank6_platform_platform1_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd34));
assign videosoc_csrbank6_platform_platform0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_platform0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd35));
assign videosoc_csrbank6_platform_target7_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target7_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd36));
assign videosoc_csrbank6_platform_target6_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target6_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd37));
assign videosoc_csrbank6_platform_target5_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target5_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd38));
assign videosoc_csrbank6_platform_target4_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target4_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd39));
assign videosoc_csrbank6_platform_target3_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target3_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd40));
assign videosoc_csrbank6_platform_target2_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target2_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd41));
assign videosoc_csrbank6_platform_target1_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd42));
assign videosoc_csrbank6_platform_target0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_platform_target0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd43));
assign videosoc_csrbank6_xadc_temperature1_r = videosoc_interface6_bank_bus_dat_w[3:0];
assign videosoc_csrbank6_xadc_temperature1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd44));
assign videosoc_csrbank6_xadc_temperature0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_xadc_temperature0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd45));
assign videosoc_csrbank6_xadc_vccint1_r = videosoc_interface6_bank_bus_dat_w[3:0];
assign videosoc_csrbank6_xadc_vccint1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd46));
assign videosoc_csrbank6_xadc_vccint0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_xadc_vccint0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd47));
assign videosoc_csrbank6_xadc_vccaux1_r = videosoc_interface6_bank_bus_dat_w[3:0];
assign videosoc_csrbank6_xadc_vccaux1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd48));
assign videosoc_csrbank6_xadc_vccaux0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_xadc_vccaux0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd49));
assign videosoc_csrbank6_xadc_vccbram1_r = videosoc_interface6_bank_bus_dat_w[3:0];
assign videosoc_csrbank6_xadc_vccbram1_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd50));
assign videosoc_csrbank6_xadc_vccbram0_r = videosoc_interface6_bank_bus_dat_w[7:0];
assign videosoc_csrbank6_xadc_vccbram0_re = ((videosoc_csrbank6_sel & videosoc_interface6_bank_bus_we) & (videosoc_interface6_bank_bus_adr[5:0] == 6'd51));
assign videosoc_csrbank6_dna_id7_w = videosoc_info_dna_status[56];
assign videosoc_csrbank6_dna_id6_w = videosoc_info_dna_status[55:48];
assign videosoc_csrbank6_dna_id5_w = videosoc_info_dna_status[47:40];
assign videosoc_csrbank6_dna_id4_w = videosoc_info_dna_status[39:32];
assign videosoc_csrbank6_dna_id3_w = videosoc_info_dna_status[31:24];
assign videosoc_csrbank6_dna_id2_w = videosoc_info_dna_status[23:16];
assign videosoc_csrbank6_dna_id1_w = videosoc_info_dna_status[15:8];
assign videosoc_csrbank6_dna_id0_w = videosoc_info_dna_status[7:0];
assign videosoc_csrbank6_git_commit19_w = videosoc_info_git_status[159:152];
assign videosoc_csrbank6_git_commit18_w = videosoc_info_git_status[151:144];
assign videosoc_csrbank6_git_commit17_w = videosoc_info_git_status[143:136];
assign videosoc_csrbank6_git_commit16_w = videosoc_info_git_status[135:128];
assign videosoc_csrbank6_git_commit15_w = videosoc_info_git_status[127:120];
assign videosoc_csrbank6_git_commit14_w = videosoc_info_git_status[119:112];
assign videosoc_csrbank6_git_commit13_w = videosoc_info_git_status[111:104];
assign videosoc_csrbank6_git_commit12_w = videosoc_info_git_status[103:96];
assign videosoc_csrbank6_git_commit11_w = videosoc_info_git_status[95:88];
assign videosoc_csrbank6_git_commit10_w = videosoc_info_git_status[87:80];
assign videosoc_csrbank6_git_commit9_w = videosoc_info_git_status[79:72];
assign videosoc_csrbank6_git_commit8_w = videosoc_info_git_status[71:64];
assign videosoc_csrbank6_git_commit7_w = videosoc_info_git_status[63:56];
assign videosoc_csrbank6_git_commit6_w = videosoc_info_git_status[55:48];
assign videosoc_csrbank6_git_commit5_w = videosoc_info_git_status[47:40];
assign videosoc_csrbank6_git_commit4_w = videosoc_info_git_status[39:32];
assign videosoc_csrbank6_git_commit3_w = videosoc_info_git_status[31:24];
assign videosoc_csrbank6_git_commit2_w = videosoc_info_git_status[23:16];
assign videosoc_csrbank6_git_commit1_w = videosoc_info_git_status[15:8];
assign videosoc_csrbank6_git_commit0_w = videosoc_info_git_status[7:0];
assign videosoc_csrbank6_platform_platform7_w = videosoc_info_platform_status[63:56];
assign videosoc_csrbank6_platform_platform6_w = videosoc_info_platform_status[55:48];
assign videosoc_csrbank6_platform_platform5_w = videosoc_info_platform_status[47:40];
assign videosoc_csrbank6_platform_platform4_w = videosoc_info_platform_status[39:32];
assign videosoc_csrbank6_platform_platform3_w = videosoc_info_platform_status[31:24];
assign videosoc_csrbank6_platform_platform2_w = videosoc_info_platform_status[23:16];
assign videosoc_csrbank6_platform_platform1_w = videosoc_info_platform_status[15:8];
assign videosoc_csrbank6_platform_platform0_w = videosoc_info_platform_status[7:0];
assign videosoc_csrbank6_platform_target7_w = videosoc_info_target_status[63:56];
assign videosoc_csrbank6_platform_target6_w = videosoc_info_target_status[55:48];
assign videosoc_csrbank6_platform_target5_w = videosoc_info_target_status[47:40];
assign videosoc_csrbank6_platform_target4_w = videosoc_info_target_status[39:32];
assign videosoc_csrbank6_platform_target3_w = videosoc_info_target_status[31:24];
assign videosoc_csrbank6_platform_target2_w = videosoc_info_target_status[23:16];
assign videosoc_csrbank6_platform_target1_w = videosoc_info_target_status[15:8];
assign videosoc_csrbank6_platform_target0_w = videosoc_info_target_status[7:0];
assign videosoc_csrbank6_xadc_temperature1_w = videosoc_info_temperature_status[11:8];
assign videosoc_csrbank6_xadc_temperature0_w = videosoc_info_temperature_status[7:0];
assign videosoc_csrbank6_xadc_vccint1_w = videosoc_info_vccint_status[11:8];
assign videosoc_csrbank6_xadc_vccint0_w = videosoc_info_vccint_status[7:0];
assign videosoc_csrbank6_xadc_vccaux1_w = videosoc_info_vccaux_status[11:8];
assign videosoc_csrbank6_xadc_vccaux0_w = videosoc_info_vccaux_status[7:0];
assign videosoc_csrbank6_xadc_vccbram1_w = videosoc_info_vccbram_status[11:8];
assign videosoc_csrbank6_xadc_vccbram0_w = videosoc_info_vccbram_status[7:0];
assign videosoc_csrbank7_sel = (videosoc_interface7_bank_bus_adr[13:9] == 4'd13);
assign videosoc_oled_spimaster_ctrl_r = videosoc_interface7_bank_bus_dat_w[0];
assign videosoc_oled_spimaster_ctrl_re = ((videosoc_csrbank7_sel & videosoc_interface7_bank_bus_we) & (videosoc_interface7_bank_bus_adr[2:0] == 1'd0));
assign videosoc_csrbank7_spi_length0_r = videosoc_interface7_bank_bus_dat_w[7:0];
assign videosoc_csrbank7_spi_length0_re = ((videosoc_csrbank7_sel & videosoc_interface7_bank_bus_we) & (videosoc_interface7_bank_bus_adr[2:0] == 1'd1));
assign videosoc_csrbank7_spi_status_r = videosoc_interface7_bank_bus_dat_w[0];
assign videosoc_csrbank7_spi_status_re = ((videosoc_csrbank7_sel & videosoc_interface7_bank_bus_we) & (videosoc_interface7_bank_bus_adr[2:0] == 2'd2));
assign videosoc_csrbank7_spi_mosi0_r = videosoc_interface7_bank_bus_dat_w[7:0];
assign videosoc_csrbank7_spi_mosi0_re = ((videosoc_csrbank7_sel & videosoc_interface7_bank_bus_we) & (videosoc_interface7_bank_bus_adr[2:0] == 2'd3));
assign videosoc_csrbank7_gpio_out0_r = videosoc_interface7_bank_bus_dat_w[3:0];
assign videosoc_csrbank7_gpio_out0_re = ((videosoc_csrbank7_sel & videosoc_interface7_bank_bus_we) & (videosoc_interface7_bank_bus_adr[2:0] == 3'd4));
assign videosoc_oled_spimaster_length_storage = videosoc_oled_spimaster_length_storage_full[7:0];
assign videosoc_csrbank7_spi_length0_w = videosoc_oled_spimaster_length_storage_full[7:0];
assign videosoc_csrbank7_spi_status_w = videosoc_oled_spimaster_status;
assign videosoc_oled_spimaster_mosi_storage = videosoc_oled_spimaster_mosi_storage_full[7:0];
assign videosoc_csrbank7_spi_mosi0_w = videosoc_oled_spimaster_mosi_storage_full[7:0];
assign videosoc_oled_storage = videosoc_oled_storage_full[3:0];
assign videosoc_csrbank7_gpio_out0_w = videosoc_oled_storage_full[3:0];
assign videosoc_csrbank8_sel = (videosoc_interface8_bank_bus_adr[13:9] == 4'd8);
assign videosoc_csrbank8_dfii_control0_r = videosoc_interface8_bank_bus_dat_w[3:0];
assign videosoc_csrbank8_dfii_control0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 1'd0));
assign videosoc_csrbank8_dfii_pi0_command0_r = videosoc_interface8_bank_bus_dat_w[5:0];
assign videosoc_csrbank8_dfii_pi0_command0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 1'd1));
assign videosoc_sdram_phaseinjector0_command_issue_r = videosoc_interface8_bank_bus_dat_w[0];
assign videosoc_sdram_phaseinjector0_command_issue_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 2'd2));
assign videosoc_csrbank8_dfii_pi0_address1_r = videosoc_interface8_bank_bus_dat_w[6:0];
assign videosoc_csrbank8_dfii_pi0_address1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 2'd3));
assign videosoc_csrbank8_dfii_pi0_address0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_address0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 3'd4));
assign videosoc_csrbank8_dfii_pi0_baddress0_r = videosoc_interface8_bank_bus_dat_w[2:0];
assign videosoc_csrbank8_dfii_pi0_baddress0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 3'd5));
assign videosoc_csrbank8_dfii_pi0_wrdata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_wrdata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 3'd6));
assign videosoc_csrbank8_dfii_pi0_wrdata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_wrdata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 3'd7));
assign videosoc_csrbank8_dfii_pi0_wrdata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_wrdata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd8));
assign videosoc_csrbank8_dfii_pi0_wrdata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_wrdata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd9));
assign videosoc_csrbank8_dfii_pi0_rddata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_rddata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd10));
assign videosoc_csrbank8_dfii_pi0_rddata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_rddata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd11));
assign videosoc_csrbank8_dfii_pi0_rddata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_rddata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd12));
assign videosoc_csrbank8_dfii_pi0_rddata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi0_rddata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd13));
assign videosoc_csrbank8_dfii_pi1_command0_r = videosoc_interface8_bank_bus_dat_w[5:0];
assign videosoc_csrbank8_dfii_pi1_command0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd14));
assign videosoc_sdram_phaseinjector1_command_issue_r = videosoc_interface8_bank_bus_dat_w[0];
assign videosoc_sdram_phaseinjector1_command_issue_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 4'd15));
assign videosoc_csrbank8_dfii_pi1_address1_r = videosoc_interface8_bank_bus_dat_w[6:0];
assign videosoc_csrbank8_dfii_pi1_address1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd16));
assign videosoc_csrbank8_dfii_pi1_address0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_address0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd17));
assign videosoc_csrbank8_dfii_pi1_baddress0_r = videosoc_interface8_bank_bus_dat_w[2:0];
assign videosoc_csrbank8_dfii_pi1_baddress0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd18));
assign videosoc_csrbank8_dfii_pi1_wrdata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_wrdata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd19));
assign videosoc_csrbank8_dfii_pi1_wrdata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_wrdata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd20));
assign videosoc_csrbank8_dfii_pi1_wrdata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_wrdata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd21));
assign videosoc_csrbank8_dfii_pi1_wrdata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_wrdata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd22));
assign videosoc_csrbank8_dfii_pi1_rddata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_rddata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd23));
assign videosoc_csrbank8_dfii_pi1_rddata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_rddata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd24));
assign videosoc_csrbank8_dfii_pi1_rddata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_rddata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd25));
assign videosoc_csrbank8_dfii_pi1_rddata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi1_rddata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd26));
assign videosoc_csrbank8_dfii_pi2_command0_r = videosoc_interface8_bank_bus_dat_w[5:0];
assign videosoc_csrbank8_dfii_pi2_command0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd27));
assign videosoc_sdram_phaseinjector2_command_issue_r = videosoc_interface8_bank_bus_dat_w[0];
assign videosoc_sdram_phaseinjector2_command_issue_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd28));
assign videosoc_csrbank8_dfii_pi2_address1_r = videosoc_interface8_bank_bus_dat_w[6:0];
assign videosoc_csrbank8_dfii_pi2_address1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd29));
assign videosoc_csrbank8_dfii_pi2_address0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_address0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd30));
assign videosoc_csrbank8_dfii_pi2_baddress0_r = videosoc_interface8_bank_bus_dat_w[2:0];
assign videosoc_csrbank8_dfii_pi2_baddress0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 5'd31));
assign videosoc_csrbank8_dfii_pi2_wrdata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_wrdata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd32));
assign videosoc_csrbank8_dfii_pi2_wrdata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_wrdata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd33));
assign videosoc_csrbank8_dfii_pi2_wrdata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_wrdata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd34));
assign videosoc_csrbank8_dfii_pi2_wrdata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_wrdata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd35));
assign videosoc_csrbank8_dfii_pi2_rddata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_rddata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd36));
assign videosoc_csrbank8_dfii_pi2_rddata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_rddata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd37));
assign videosoc_csrbank8_dfii_pi2_rddata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_rddata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd38));
assign videosoc_csrbank8_dfii_pi2_rddata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi2_rddata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd39));
assign videosoc_csrbank8_dfii_pi3_command0_r = videosoc_interface8_bank_bus_dat_w[5:0];
assign videosoc_csrbank8_dfii_pi3_command0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd40));
assign videosoc_sdram_phaseinjector3_command_issue_r = videosoc_interface8_bank_bus_dat_w[0];
assign videosoc_sdram_phaseinjector3_command_issue_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd41));
assign videosoc_csrbank8_dfii_pi3_address1_r = videosoc_interface8_bank_bus_dat_w[6:0];
assign videosoc_csrbank8_dfii_pi3_address1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd42));
assign videosoc_csrbank8_dfii_pi3_address0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_address0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd43));
assign videosoc_csrbank8_dfii_pi3_baddress0_r = videosoc_interface8_bank_bus_dat_w[2:0];
assign videosoc_csrbank8_dfii_pi3_baddress0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd44));
assign videosoc_csrbank8_dfii_pi3_wrdata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_wrdata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd45));
assign videosoc_csrbank8_dfii_pi3_wrdata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_wrdata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd46));
assign videosoc_csrbank8_dfii_pi3_wrdata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_wrdata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd47));
assign videosoc_csrbank8_dfii_pi3_wrdata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_wrdata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd48));
assign videosoc_csrbank8_dfii_pi3_rddata3_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_rddata3_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd49));
assign videosoc_csrbank8_dfii_pi3_rddata2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_rddata2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd50));
assign videosoc_csrbank8_dfii_pi3_rddata1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_rddata1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd51));
assign videosoc_csrbank8_dfii_pi3_rddata0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_dfii_pi3_rddata0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd52));
assign videosoc_sdram_bandwidth_update_r = videosoc_interface8_bank_bus_dat_w[0];
assign videosoc_sdram_bandwidth_update_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd53));
assign videosoc_csrbank8_controller_bandwidth_nreads2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_controller_bandwidth_nreads2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd54));
assign videosoc_csrbank8_controller_bandwidth_nreads1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_controller_bandwidth_nreads1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd55));
assign videosoc_csrbank8_controller_bandwidth_nreads0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_controller_bandwidth_nreads0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd56));
assign videosoc_csrbank8_controller_bandwidth_nwrites2_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_controller_bandwidth_nwrites2_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd57));
assign videosoc_csrbank8_controller_bandwidth_nwrites1_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_controller_bandwidth_nwrites1_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd58));
assign videosoc_csrbank8_controller_bandwidth_nwrites0_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_controller_bandwidth_nwrites0_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd59));
assign videosoc_csrbank8_controller_bandwidth_data_width_r = videosoc_interface8_bank_bus_dat_w[7:0];
assign videosoc_csrbank8_controller_bandwidth_data_width_re = ((videosoc_csrbank8_sel & videosoc_interface8_bank_bus_we) & (videosoc_interface8_bank_bus_adr[5:0] == 6'd60));
assign videosoc_sdram_storage = videosoc_sdram_storage_full[3:0];
assign videosoc_csrbank8_dfii_control0_w = videosoc_sdram_storage_full[3:0];
assign videosoc_sdram_phaseinjector0_command_storage = videosoc_sdram_phaseinjector0_command_storage_full[5:0];
assign videosoc_csrbank8_dfii_pi0_command0_w = videosoc_sdram_phaseinjector0_command_storage_full[5:0];
assign videosoc_sdram_phaseinjector0_address_storage = videosoc_sdram_phaseinjector0_address_storage_full[14:0];
assign videosoc_csrbank8_dfii_pi0_address1_w = videosoc_sdram_phaseinjector0_address_storage_full[14:8];
assign videosoc_csrbank8_dfii_pi0_address0_w = videosoc_sdram_phaseinjector0_address_storage_full[7:0];
assign videosoc_sdram_phaseinjector0_baddress_storage = videosoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign videosoc_csrbank8_dfii_pi0_baddress0_w = videosoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign videosoc_sdram_phaseinjector0_wrdata_storage = videosoc_sdram_phaseinjector0_wrdata_storage_full[31:0];
assign videosoc_csrbank8_dfii_pi0_wrdata3_w = videosoc_sdram_phaseinjector0_wrdata_storage_full[31:24];
assign videosoc_csrbank8_dfii_pi0_wrdata2_w = videosoc_sdram_phaseinjector0_wrdata_storage_full[23:16];
assign videosoc_csrbank8_dfii_pi0_wrdata1_w = videosoc_sdram_phaseinjector0_wrdata_storage_full[15:8];
assign videosoc_csrbank8_dfii_pi0_wrdata0_w = videosoc_sdram_phaseinjector0_wrdata_storage_full[7:0];
assign videosoc_csrbank8_dfii_pi0_rddata3_w = videosoc_sdram_phaseinjector0_status[31:24];
assign videosoc_csrbank8_dfii_pi0_rddata2_w = videosoc_sdram_phaseinjector0_status[23:16];
assign videosoc_csrbank8_dfii_pi0_rddata1_w = videosoc_sdram_phaseinjector0_status[15:8];
assign videosoc_csrbank8_dfii_pi0_rddata0_w = videosoc_sdram_phaseinjector0_status[7:0];
assign videosoc_sdram_phaseinjector1_command_storage = videosoc_sdram_phaseinjector1_command_storage_full[5:0];
assign videosoc_csrbank8_dfii_pi1_command0_w = videosoc_sdram_phaseinjector1_command_storage_full[5:0];
assign videosoc_sdram_phaseinjector1_address_storage = videosoc_sdram_phaseinjector1_address_storage_full[14:0];
assign videosoc_csrbank8_dfii_pi1_address1_w = videosoc_sdram_phaseinjector1_address_storage_full[14:8];
assign videosoc_csrbank8_dfii_pi1_address0_w = videosoc_sdram_phaseinjector1_address_storage_full[7:0];
assign videosoc_sdram_phaseinjector1_baddress_storage = videosoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign videosoc_csrbank8_dfii_pi1_baddress0_w = videosoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign videosoc_sdram_phaseinjector1_wrdata_storage = videosoc_sdram_phaseinjector1_wrdata_storage_full[31:0];
assign videosoc_csrbank8_dfii_pi1_wrdata3_w = videosoc_sdram_phaseinjector1_wrdata_storage_full[31:24];
assign videosoc_csrbank8_dfii_pi1_wrdata2_w = videosoc_sdram_phaseinjector1_wrdata_storage_full[23:16];
assign videosoc_csrbank8_dfii_pi1_wrdata1_w = videosoc_sdram_phaseinjector1_wrdata_storage_full[15:8];
assign videosoc_csrbank8_dfii_pi1_wrdata0_w = videosoc_sdram_phaseinjector1_wrdata_storage_full[7:0];
assign videosoc_csrbank8_dfii_pi1_rddata3_w = videosoc_sdram_phaseinjector1_status[31:24];
assign videosoc_csrbank8_dfii_pi1_rddata2_w = videosoc_sdram_phaseinjector1_status[23:16];
assign videosoc_csrbank8_dfii_pi1_rddata1_w = videosoc_sdram_phaseinjector1_status[15:8];
assign videosoc_csrbank8_dfii_pi1_rddata0_w = videosoc_sdram_phaseinjector1_status[7:0];
assign videosoc_sdram_phaseinjector2_command_storage = videosoc_sdram_phaseinjector2_command_storage_full[5:0];
assign videosoc_csrbank8_dfii_pi2_command0_w = videosoc_sdram_phaseinjector2_command_storage_full[5:0];
assign videosoc_sdram_phaseinjector2_address_storage = videosoc_sdram_phaseinjector2_address_storage_full[14:0];
assign videosoc_csrbank8_dfii_pi2_address1_w = videosoc_sdram_phaseinjector2_address_storage_full[14:8];
assign videosoc_csrbank8_dfii_pi2_address0_w = videosoc_sdram_phaseinjector2_address_storage_full[7:0];
assign videosoc_sdram_phaseinjector2_baddress_storage = videosoc_sdram_phaseinjector2_baddress_storage_full[2:0];
assign videosoc_csrbank8_dfii_pi2_baddress0_w = videosoc_sdram_phaseinjector2_baddress_storage_full[2:0];
assign videosoc_sdram_phaseinjector2_wrdata_storage = videosoc_sdram_phaseinjector2_wrdata_storage_full[31:0];
assign videosoc_csrbank8_dfii_pi2_wrdata3_w = videosoc_sdram_phaseinjector2_wrdata_storage_full[31:24];
assign videosoc_csrbank8_dfii_pi2_wrdata2_w = videosoc_sdram_phaseinjector2_wrdata_storage_full[23:16];
assign videosoc_csrbank8_dfii_pi2_wrdata1_w = videosoc_sdram_phaseinjector2_wrdata_storage_full[15:8];
assign videosoc_csrbank8_dfii_pi2_wrdata0_w = videosoc_sdram_phaseinjector2_wrdata_storage_full[7:0];
assign videosoc_csrbank8_dfii_pi2_rddata3_w = videosoc_sdram_phaseinjector2_status[31:24];
assign videosoc_csrbank8_dfii_pi2_rddata2_w = videosoc_sdram_phaseinjector2_status[23:16];
assign videosoc_csrbank8_dfii_pi2_rddata1_w = videosoc_sdram_phaseinjector2_status[15:8];
assign videosoc_csrbank8_dfii_pi2_rddata0_w = videosoc_sdram_phaseinjector2_status[7:0];
assign videosoc_sdram_phaseinjector3_command_storage = videosoc_sdram_phaseinjector3_command_storage_full[5:0];
assign videosoc_csrbank8_dfii_pi3_command0_w = videosoc_sdram_phaseinjector3_command_storage_full[5:0];
assign videosoc_sdram_phaseinjector3_address_storage = videosoc_sdram_phaseinjector3_address_storage_full[14:0];
assign videosoc_csrbank8_dfii_pi3_address1_w = videosoc_sdram_phaseinjector3_address_storage_full[14:8];
assign videosoc_csrbank8_dfii_pi3_address0_w = videosoc_sdram_phaseinjector3_address_storage_full[7:0];
assign videosoc_sdram_phaseinjector3_baddress_storage = videosoc_sdram_phaseinjector3_baddress_storage_full[2:0];
assign videosoc_csrbank8_dfii_pi3_baddress0_w = videosoc_sdram_phaseinjector3_baddress_storage_full[2:0];
assign videosoc_sdram_phaseinjector3_wrdata_storage = videosoc_sdram_phaseinjector3_wrdata_storage_full[31:0];
assign videosoc_csrbank8_dfii_pi3_wrdata3_w = videosoc_sdram_phaseinjector3_wrdata_storage_full[31:24];
assign videosoc_csrbank8_dfii_pi3_wrdata2_w = videosoc_sdram_phaseinjector3_wrdata_storage_full[23:16];
assign videosoc_csrbank8_dfii_pi3_wrdata1_w = videosoc_sdram_phaseinjector3_wrdata_storage_full[15:8];
assign videosoc_csrbank8_dfii_pi3_wrdata0_w = videosoc_sdram_phaseinjector3_wrdata_storage_full[7:0];
assign videosoc_csrbank8_dfii_pi3_rddata3_w = videosoc_sdram_phaseinjector3_status[31:24];
assign videosoc_csrbank8_dfii_pi3_rddata2_w = videosoc_sdram_phaseinjector3_status[23:16];
assign videosoc_csrbank8_dfii_pi3_rddata1_w = videosoc_sdram_phaseinjector3_status[15:8];
assign videosoc_csrbank8_dfii_pi3_rddata0_w = videosoc_sdram_phaseinjector3_status[7:0];
assign videosoc_csrbank8_controller_bandwidth_nreads2_w = videosoc_sdram_bandwidth_nreads_status[23:16];
assign videosoc_csrbank8_controller_bandwidth_nreads1_w = videosoc_sdram_bandwidth_nreads_status[15:8];
assign videosoc_csrbank8_controller_bandwidth_nreads0_w = videosoc_sdram_bandwidth_nreads_status[7:0];
assign videosoc_csrbank8_controller_bandwidth_nwrites2_w = videosoc_sdram_bandwidth_nwrites_status[23:16];
assign videosoc_csrbank8_controller_bandwidth_nwrites1_w = videosoc_sdram_bandwidth_nwrites_status[15:8];
assign videosoc_csrbank8_controller_bandwidth_nwrites0_w = videosoc_sdram_bandwidth_nwrites_status[7:0];
assign videosoc_csrbank8_controller_bandwidth_data_width_w = videosoc_sdram_bandwidth_data_width_status[7:0];
assign videosoc_csrbank9_sel = (videosoc_interface9_bank_bus_adr[13:9] == 4'd10);
assign videosoc_csrbank9_bitbang0_r = videosoc_interface9_bank_bus_dat_w[3:0];
assign videosoc_csrbank9_bitbang0_re = ((videosoc_csrbank9_sel & videosoc_interface9_bank_bus_we) & (videosoc_interface9_bank_bus_adr[1:0] == 1'd0));
assign videosoc_csrbank9_miso_r = videosoc_interface9_bank_bus_dat_w[0];
assign videosoc_csrbank9_miso_re = ((videosoc_csrbank9_sel & videosoc_interface9_bank_bus_we) & (videosoc_interface9_bank_bus_adr[1:0] == 1'd1));
assign videosoc_csrbank9_bitbang_en0_r = videosoc_interface9_bank_bus_dat_w[0];
assign videosoc_csrbank9_bitbang_en0_re = ((videosoc_csrbank9_sel & videosoc_interface9_bank_bus_we) & (videosoc_interface9_bank_bus_adr[1:0] == 2'd2));
assign videosoc_bitbang_storage = videosoc_bitbang_storage_full[3:0];
assign videosoc_csrbank9_bitbang0_w = videosoc_bitbang_storage_full[3:0];
assign videosoc_csrbank9_miso_w = videosoc_miso_status;
assign videosoc_bitbang_en_storage = videosoc_bitbang_en_storage_full;
assign videosoc_csrbank9_bitbang_en0_w = videosoc_bitbang_en_storage_full;
assign videosoc_csrbank10_sel = (videosoc_interface10_bank_bus_adr[13:9] == 3'd4);
assign videosoc_csrbank10_load3_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_load3_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 1'd0));
assign videosoc_csrbank10_load2_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_load2_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 1'd1));
assign videosoc_csrbank10_load1_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_load1_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 2'd2));
assign videosoc_csrbank10_load0_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_load0_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 2'd3));
assign videosoc_csrbank10_reload3_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_reload3_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 3'd4));
assign videosoc_csrbank10_reload2_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_reload2_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 3'd5));
assign videosoc_csrbank10_reload1_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_reload1_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 3'd6));
assign videosoc_csrbank10_reload0_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_reload0_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 3'd7));
assign videosoc_csrbank10_en0_r = videosoc_interface10_bank_bus_dat_w[0];
assign videosoc_csrbank10_en0_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd8));
assign videosoc_videosoc_update_value_r = videosoc_interface10_bank_bus_dat_w[0];
assign videosoc_videosoc_update_value_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd9));
assign videosoc_csrbank10_value3_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_value3_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd10));
assign videosoc_csrbank10_value2_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_value2_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd11));
assign videosoc_csrbank10_value1_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_value1_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd12));
assign videosoc_csrbank10_value0_r = videosoc_interface10_bank_bus_dat_w[7:0];
assign videosoc_csrbank10_value0_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd13));
assign videosoc_videosoc_eventmanager_status_r = videosoc_interface10_bank_bus_dat_w[0];
assign videosoc_videosoc_eventmanager_status_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd14));
assign videosoc_videosoc_eventmanager_pending_r = videosoc_interface10_bank_bus_dat_w[0];
assign videosoc_videosoc_eventmanager_pending_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 4'd15));
assign videosoc_csrbank10_ev_enable0_r = videosoc_interface10_bank_bus_dat_w[0];
assign videosoc_csrbank10_ev_enable0_re = ((videosoc_csrbank10_sel & videosoc_interface10_bank_bus_we) & (videosoc_interface10_bank_bus_adr[4:0] == 5'd16));
assign videosoc_videosoc_load_storage = videosoc_videosoc_load_storage_full[31:0];
assign videosoc_csrbank10_load3_w = videosoc_videosoc_load_storage_full[31:24];
assign videosoc_csrbank10_load2_w = videosoc_videosoc_load_storage_full[23:16];
assign videosoc_csrbank10_load1_w = videosoc_videosoc_load_storage_full[15:8];
assign videosoc_csrbank10_load0_w = videosoc_videosoc_load_storage_full[7:0];
assign videosoc_videosoc_reload_storage = videosoc_videosoc_reload_storage_full[31:0];
assign videosoc_csrbank10_reload3_w = videosoc_videosoc_reload_storage_full[31:24];
assign videosoc_csrbank10_reload2_w = videosoc_videosoc_reload_storage_full[23:16];
assign videosoc_csrbank10_reload1_w = videosoc_videosoc_reload_storage_full[15:8];
assign videosoc_csrbank10_reload0_w = videosoc_videosoc_reload_storage_full[7:0];
assign videosoc_videosoc_en_storage = videosoc_videosoc_en_storage_full;
assign videosoc_csrbank10_en0_w = videosoc_videosoc_en_storage_full;
assign videosoc_csrbank10_value3_w = videosoc_videosoc_value_status[31:24];
assign videosoc_csrbank10_value2_w = videosoc_videosoc_value_status[23:16];
assign videosoc_csrbank10_value1_w = videosoc_videosoc_value_status[15:8];
assign videosoc_csrbank10_value0_w = videosoc_videosoc_value_status[7:0];
assign videosoc_videosoc_eventmanager_storage = videosoc_videosoc_eventmanager_storage_full;
assign videosoc_csrbank10_ev_enable0_w = videosoc_videosoc_eventmanager_storage_full;
assign videosoc_csrbank11_sel = (videosoc_interface11_bank_bus_adr[13:9] == 2'd2);
assign videosoc_uart_rxtx_r = videosoc_interface11_bank_bus_dat_w[7:0];
assign videosoc_uart_rxtx_re = ((videosoc_csrbank11_sel & videosoc_interface11_bank_bus_we) & (videosoc_interface11_bank_bus_adr[2:0] == 1'd0));
assign videosoc_csrbank11_txfull_r = videosoc_interface11_bank_bus_dat_w[0];
assign videosoc_csrbank11_txfull_re = ((videosoc_csrbank11_sel & videosoc_interface11_bank_bus_we) & (videosoc_interface11_bank_bus_adr[2:0] == 1'd1));
assign videosoc_csrbank11_rxempty_r = videosoc_interface11_bank_bus_dat_w[0];
assign videosoc_csrbank11_rxempty_re = ((videosoc_csrbank11_sel & videosoc_interface11_bank_bus_we) & (videosoc_interface11_bank_bus_adr[2:0] == 2'd2));
assign videosoc_uart_status_r = videosoc_interface11_bank_bus_dat_w[1:0];
assign videosoc_uart_status_re = ((videosoc_csrbank11_sel & videosoc_interface11_bank_bus_we) & (videosoc_interface11_bank_bus_adr[2:0] == 2'd3));
assign videosoc_uart_pending_r = videosoc_interface11_bank_bus_dat_w[1:0];
assign videosoc_uart_pending_re = ((videosoc_csrbank11_sel & videosoc_interface11_bank_bus_we) & (videosoc_interface11_bank_bus_adr[2:0] == 3'd4));
assign videosoc_csrbank11_ev_enable0_r = videosoc_interface11_bank_bus_dat_w[1:0];
assign videosoc_csrbank11_ev_enable0_re = ((videosoc_csrbank11_sel & videosoc_interface11_bank_bus_we) & (videosoc_interface11_bank_bus_adr[2:0] == 3'd5));
assign videosoc_csrbank11_txfull_w = videosoc_uart_txfull_status;
assign videosoc_csrbank11_rxempty_w = videosoc_uart_rxempty_status;
assign videosoc_uart_storage = videosoc_uart_storage_full[1:0];
assign videosoc_csrbank11_ev_enable0_w = videosoc_uart_storage_full[1:0];
assign videosoc_csrbank12_sel = (videosoc_interface12_bank_bus_adr[13:9] == 1'd1);
assign videosoc_csrbank12_tuning_word3_r = videosoc_interface12_bank_bus_dat_w[7:0];
assign videosoc_csrbank12_tuning_word3_re = ((videosoc_csrbank12_sel & videosoc_interface12_bank_bus_we) & (videosoc_interface12_bank_bus_adr[1:0] == 1'd0));
assign videosoc_csrbank12_tuning_word2_r = videosoc_interface12_bank_bus_dat_w[7:0];
assign videosoc_csrbank12_tuning_word2_re = ((videosoc_csrbank12_sel & videosoc_interface12_bank_bus_we) & (videosoc_interface12_bank_bus_adr[1:0] == 1'd1));
assign videosoc_csrbank12_tuning_word1_r = videosoc_interface12_bank_bus_dat_w[7:0];
assign videosoc_csrbank12_tuning_word1_re = ((videosoc_csrbank12_sel & videosoc_interface12_bank_bus_we) & (videosoc_interface12_bank_bus_adr[1:0] == 2'd2));
assign videosoc_csrbank12_tuning_word0_r = videosoc_interface12_bank_bus_dat_w[7:0];
assign videosoc_csrbank12_tuning_word0_re = ((videosoc_csrbank12_sel & videosoc_interface12_bank_bus_we) & (videosoc_interface12_bank_bus_adr[1:0] == 2'd3));
assign videosoc_uart_phy_storage = videosoc_uart_phy_storage_full[31:0];
assign videosoc_csrbank12_tuning_word3_w = videosoc_uart_phy_storage_full[31:24];
assign videosoc_csrbank12_tuning_word2_w = videosoc_uart_phy_storage_full[23:16];
assign videosoc_csrbank12_tuning_word1_w = videosoc_uart_phy_storage_full[15:8];
assign videosoc_csrbank12_tuning_word0_w = videosoc_uart_phy_storage_full[7:0];
assign videosoc_interface0_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface1_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface2_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface3_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface4_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface5_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface6_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface7_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface8_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface9_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface10_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface11_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface12_bank_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface0_sram_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface1_sram_bus_adr = videosoc_videosoc_interface_adr;
assign videosoc_interface0_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface1_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface2_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface3_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface4_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface5_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface6_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface7_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface8_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface9_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface10_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface11_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface12_bank_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface0_sram_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface1_sram_bus_we = videosoc_videosoc_interface_we;
assign videosoc_interface0_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface1_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface2_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface3_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface4_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface5_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface6_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface7_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface8_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface9_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface10_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface11_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface12_bank_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface0_sram_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_interface1_sram_bus_dat_w = videosoc_videosoc_interface_dat_w;
assign videosoc_videosoc_interface_dat_r = ((((((((((((((videosoc_interface0_bank_bus_dat_r | videosoc_interface1_bank_bus_dat_r) | videosoc_interface2_bank_bus_dat_r) | videosoc_interface3_bank_bus_dat_r) | videosoc_interface4_bank_bus_dat_r) | videosoc_interface5_bank_bus_dat_r) | videosoc_interface6_bank_bus_dat_r) | videosoc_interface7_bank_bus_dat_r) | videosoc_interface8_bank_bus_dat_r) | videosoc_interface9_bank_bus_dat_r) | videosoc_interface10_bank_bus_dat_r) | videosoc_interface11_bank_bus_dat_r) | videosoc_interface12_bank_bus_dat_r) | videosoc_interface0_sram_bus_dat_r) | videosoc_interface1_sram_bus_dat_r);
always @(*) begin
	comb_rhs_array_muxed0 <= 1'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[0];
		end
		1'd1: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[1];
		end
		2'd2: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[2];
		end
		2'd3: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[3];
		end
		3'd4: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[4];
		end
		3'd5: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[5];
		end
		3'd6: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[6];
		end
		default: begin
			comb_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_valids[7];
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed1 <= 15'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			comb_rhs_array_muxed1 <= videosoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed2 <= 3'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			comb_rhs_array_muxed2 <= videosoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed3 <= 1'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			comb_rhs_array_muxed3 <= videosoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed4 <= 1'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			comb_rhs_array_muxed4 <= videosoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed5 <= 1'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			comb_rhs_array_muxed5 <= videosoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	comb_t_array_muxed0 <= 1'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			comb_t_array_muxed0 <= videosoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	comb_t_array_muxed1 <= 1'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			comb_t_array_muxed1 <= videosoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	comb_t_array_muxed2 <= 1'd0;
	case (videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			comb_t_array_muxed2 <= videosoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed6 <= 1'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[0];
		end
		1'd1: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[1];
		end
		2'd2: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[2];
		end
		2'd3: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[3];
		end
		3'd4: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[4];
		end
		3'd5: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[5];
		end
		3'd6: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[6];
		end
		default: begin
			comb_rhs_array_muxed6 <= videosoc_sdram_choose_req_valids[7];
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed7 <= 15'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			comb_rhs_array_muxed7 <= videosoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed8 <= 3'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			comb_rhs_array_muxed8 <= videosoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed9 <= 1'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			comb_rhs_array_muxed9 <= videosoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed10 <= 1'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			comb_rhs_array_muxed10 <= videosoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed11 <= 1'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			comb_rhs_array_muxed11 <= videosoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	comb_t_array_muxed3 <= 1'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			comb_t_array_muxed3 <= videosoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	comb_t_array_muxed4 <= 1'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			comb_t_array_muxed4 <= videosoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	comb_t_array_muxed5 <= 1'd0;
	case (videosoc_sdram_choose_req_grant)
		1'd0: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			comb_t_array_muxed5 <= videosoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed12 <= 22'd0;
	case (roundrobin0_grant)
		1'd0: begin
			comb_rhs_array_muxed12 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed12 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed12 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed13 <= 1'd0;
	case (roundrobin0_grant)
		1'd0: begin
			comb_rhs_array_muxed13 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed13 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed13 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed14 <= 1'd0;
	case (roundrobin0_grant)
		1'd0: begin
			comb_rhs_array_muxed14 <= (((cba0 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed14 <= (((cba1 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed14 <= (((cba2 == 1'd0) & (~(((((((1'd0 | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed15 <= 22'd0;
	case (roundrobin1_grant)
		1'd0: begin
			comb_rhs_array_muxed15 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed15 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed15 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed16 <= 1'd0;
	case (roundrobin1_grant)
		1'd0: begin
			comb_rhs_array_muxed16 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed16 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed16 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed17 <= 1'd0;
	case (roundrobin1_grant)
		1'd0: begin
			comb_rhs_array_muxed17 <= (((cba0 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed17 <= (((cba1 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed17 <= (((cba2 == 1'd1) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed18 <= 22'd0;
	case (roundrobin2_grant)
		1'd0: begin
			comb_rhs_array_muxed18 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed18 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed18 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed19 <= 1'd0;
	case (roundrobin2_grant)
		1'd0: begin
			comb_rhs_array_muxed19 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed19 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed19 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed20 <= 1'd0;
	case (roundrobin2_grant)
		1'd0: begin
			comb_rhs_array_muxed20 <= (((cba0 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed20 <= (((cba1 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed20 <= (((cba2 == 2'd2) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed21 <= 22'd0;
	case (roundrobin3_grant)
		1'd0: begin
			comb_rhs_array_muxed21 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed21 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed21 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed22 <= 1'd0;
	case (roundrobin3_grant)
		1'd0: begin
			comb_rhs_array_muxed22 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed22 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed22 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed23 <= 1'd0;
	case (roundrobin3_grant)
		1'd0: begin
			comb_rhs_array_muxed23 <= (((cba0 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed23 <= (((cba1 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed23 <= (((cba2 == 2'd3) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed24 <= 22'd0;
	case (roundrobin4_grant)
		1'd0: begin
			comb_rhs_array_muxed24 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed24 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed24 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed25 <= 1'd0;
	case (roundrobin4_grant)
		1'd0: begin
			comb_rhs_array_muxed25 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed25 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed25 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed26 <= 1'd0;
	case (roundrobin4_grant)
		1'd0: begin
			comb_rhs_array_muxed26 <= (((cba0 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed26 <= (((cba1 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed26 <= (((cba2 == 3'd4) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed27 <= 22'd0;
	case (roundrobin5_grant)
		1'd0: begin
			comb_rhs_array_muxed27 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed27 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed27 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed28 <= 1'd0;
	case (roundrobin5_grant)
		1'd0: begin
			comb_rhs_array_muxed28 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed28 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed28 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed29 <= 1'd0;
	case (roundrobin5_grant)
		1'd0: begin
			comb_rhs_array_muxed29 <= (((cba0 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed29 <= (((cba1 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed29 <= (((cba2 == 3'd5) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed30 <= 22'd0;
	case (roundrobin6_grant)
		1'd0: begin
			comb_rhs_array_muxed30 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed30 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed30 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed31 <= 1'd0;
	case (roundrobin6_grant)
		1'd0: begin
			comb_rhs_array_muxed31 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed31 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed31 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed32 <= 1'd0;
	case (roundrobin6_grant)
		1'd0: begin
			comb_rhs_array_muxed32 <= (((cba0 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed32 <= (((cba1 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed32 <= (((cba2 == 3'd6) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank7_lock & (roundrobin7_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed33 <= 22'd0;
	case (roundrobin7_grant)
		1'd0: begin
			comb_rhs_array_muxed33 <= rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed33 <= rca1;
		end
		default: begin
			comb_rhs_array_muxed33 <= rca2;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed34 <= 1'd0;
	case (roundrobin7_grant)
		1'd0: begin
			comb_rhs_array_muxed34 <= videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed34 <= litedramcrossbar_cmd_payload_we;
		end
		default: begin
			comb_rhs_array_muxed34 <= hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed35 <= 1'd0;
	case (roundrobin7_grant)
		1'd0: begin
			comb_rhs_array_muxed35 <= (((cba0 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd0))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd0))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd0))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd0))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd0))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd0))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd0))))) & videosoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed35 <= (((cba1 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 1'd1))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 1'd1))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 1'd1))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 1'd1))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 1'd1))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 1'd1))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 1'd1))))) & litedramcrossbar_cmd_valid);
		end
		default: begin
			comb_rhs_array_muxed35 <= (((cba2 == 3'd7) & (~(((((((1'd0 | (videosoc_sdram_interface_bank0_lock & (roundrobin0_grant == 2'd2))) | (videosoc_sdram_interface_bank1_lock & (roundrobin1_grant == 2'd2))) | (videosoc_sdram_interface_bank2_lock & (roundrobin2_grant == 2'd2))) | (videosoc_sdram_interface_bank3_lock & (roundrobin3_grant == 2'd2))) | (videosoc_sdram_interface_bank4_lock & (roundrobin4_grant == 2'd2))) | (videosoc_sdram_interface_bank5_lock & (roundrobin5_grant == 2'd2))) | (videosoc_sdram_interface_bank6_lock & (roundrobin6_grant == 2'd2))))) & hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed36 <= 25'd0;
	case (dma_slot_array_current_slot)
		1'd0: begin
			comb_rhs_array_muxed36 <= dma_slot_array_slot0_address;
		end
		default: begin
			comb_rhs_array_muxed36 <= dma_slot_array_slot1_address;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed37 <= 1'd0;
	case (dma_slot_array_current_slot)
		1'd0: begin
			comb_rhs_array_muxed37 <= dma_slot_array_slot0_address_valid;
		end
		default: begin
			comb_rhs_array_muxed37 <= dma_slot_array_slot1_address_valid;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed38 <= 30'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed38 <= videosoc_interface1_wb_sdram_adr;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed39 <= 32'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed39 <= videosoc_interface1_wb_sdram_dat_w;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed40 <= 4'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed40 <= videosoc_interface1_wb_sdram_sel;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed41 <= 1'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed41 <= videosoc_interface1_wb_sdram_cyc;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed42 <= 1'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed42 <= videosoc_interface1_wb_sdram_stb;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed43 <= 1'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed43 <= videosoc_interface1_wb_sdram_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed44 <= 3'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed44 <= videosoc_interface1_wb_sdram_cti;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed45 <= 2'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed45 <= videosoc_interface1_wb_sdram_bte;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed46 <= 30'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed46 <= videosoc_videosoc_ibus_adr;
		end
		1'd1: begin
			comb_rhs_array_muxed46 <= videosoc_videosoc_dbus_adr;
		end
		default: begin
			comb_rhs_array_muxed46 <= videosoc_bridge_wishbone_adr;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed47 <= 32'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed47 <= videosoc_videosoc_ibus_dat_w;
		end
		1'd1: begin
			comb_rhs_array_muxed47 <= videosoc_videosoc_dbus_dat_w;
		end
		default: begin
			comb_rhs_array_muxed47 <= videosoc_bridge_wishbone_dat_w;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed48 <= 4'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed48 <= videosoc_videosoc_ibus_sel;
		end
		1'd1: begin
			comb_rhs_array_muxed48 <= videosoc_videosoc_dbus_sel;
		end
		default: begin
			comb_rhs_array_muxed48 <= videosoc_bridge_wishbone_sel;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed49 <= 1'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed49 <= videosoc_videosoc_ibus_cyc;
		end
		1'd1: begin
			comb_rhs_array_muxed49 <= videosoc_videosoc_dbus_cyc;
		end
		default: begin
			comb_rhs_array_muxed49 <= videosoc_bridge_wishbone_cyc;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed50 <= 1'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed50 <= videosoc_videosoc_ibus_stb;
		end
		1'd1: begin
			comb_rhs_array_muxed50 <= videosoc_videosoc_dbus_stb;
		end
		default: begin
			comb_rhs_array_muxed50 <= videosoc_bridge_wishbone_stb;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed51 <= 1'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed51 <= videosoc_videosoc_ibus_we;
		end
		1'd1: begin
			comb_rhs_array_muxed51 <= videosoc_videosoc_dbus_we;
		end
		default: begin
			comb_rhs_array_muxed51 <= videosoc_bridge_wishbone_we;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed52 <= 3'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed52 <= videosoc_videosoc_ibus_cti;
		end
		1'd1: begin
			comb_rhs_array_muxed52 <= videosoc_videosoc_dbus_cti;
		end
		default: begin
			comb_rhs_array_muxed52 <= videosoc_bridge_wishbone_cti;
		end
	endcase
end
always @(*) begin
	comb_rhs_array_muxed53 <= 2'd0;
	case (videosoc_grant)
		1'd0: begin
			comb_rhs_array_muxed53 <= videosoc_videosoc_ibus_bte;
		end
		1'd1: begin
			comb_rhs_array_muxed53 <= videosoc_videosoc_dbus_bte;
		end
		default: begin
			comb_rhs_array_muxed53 <= videosoc_bridge_wishbone_bte;
		end
	endcase
end
always @(*) begin
	sync_f_array_muxed0 <= 10'd0;
	case (hdmi_out0_driver_hdmi_phy_es0_new_c2)
		1'd0: begin
			sync_f_array_muxed0 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed0 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed0 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed0 <= 10'd683;
		end
	endcase
end
always @(*) begin
	sync_f_array_muxed1 <= 10'd0;
	case (hdmi_out0_driver_hdmi_phy_es1_new_c2)
		1'd0: begin
			sync_f_array_muxed1 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed1 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed1 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed1 <= 10'd683;
		end
	endcase
end
always @(*) begin
	sync_f_array_muxed2 <= 10'd0;
	case (hdmi_out0_driver_hdmi_phy_es2_new_c2)
		1'd0: begin
			sync_f_array_muxed2 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed2 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed2 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed2 <= 10'd683;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed0 <= 15'd0;
	case (videosoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed0 <= videosoc_sdram_nop_a;
		end
		1'd1: begin
			sync_rhs_array_muxed0 <= videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			sync_rhs_array_muxed0 <= videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			sync_rhs_array_muxed0 <= videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed1 <= 3'd0;
	case (videosoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed1 <= videosoc_sdram_nop_ba;
		end
		1'd1: begin
			sync_rhs_array_muxed1 <= videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			sync_rhs_array_muxed1 <= videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			sync_rhs_array_muxed1 <= videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed2 <= 1'd0;
	case (videosoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed2 <= videosoc_sdram_nop_cas;
		end
		1'd1: begin
			sync_rhs_array_muxed2 <= videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			sync_rhs_array_muxed2 <= videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			sync_rhs_array_muxed2 <= videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed3 <= 1'd0;
	case (videosoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed3 <= videosoc_sdram_nop_ras;
		end
		1'd1: begin
			sync_rhs_array_muxed3 <= videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			sync_rhs_array_muxed3 <= videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			sync_rhs_array_muxed3 <= videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed4 <= 1'd0;
	case (videosoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed4 <= videosoc_sdram_nop_we;
		end
		1'd1: begin
			sync_rhs_array_muxed4 <= videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			sync_rhs_array_muxed4 <= videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			sync_rhs_array_muxed4 <= videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed5 <= 1'd0;
	case (videosoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed5 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed5 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			sync_rhs_array_muxed5 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			sync_rhs_array_muxed5 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed6 <= 1'd0;
	case (videosoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed6 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed6 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			sync_rhs_array_muxed6 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			sync_rhs_array_muxed6 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed7 <= 15'd0;
	case (videosoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed7 <= videosoc_sdram_nop_a;
		end
		1'd1: begin
			sync_rhs_array_muxed7 <= videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			sync_rhs_array_muxed7 <= videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			sync_rhs_array_muxed7 <= videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed8 <= 3'd0;
	case (videosoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed8 <= videosoc_sdram_nop_ba;
		end
		1'd1: begin
			sync_rhs_array_muxed8 <= videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			sync_rhs_array_muxed8 <= videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			sync_rhs_array_muxed8 <= videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed9 <= 1'd0;
	case (videosoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed9 <= videosoc_sdram_nop_cas;
		end
		1'd1: begin
			sync_rhs_array_muxed9 <= videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			sync_rhs_array_muxed9 <= videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			sync_rhs_array_muxed9 <= videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed10 <= 1'd0;
	case (videosoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed10 <= videosoc_sdram_nop_ras;
		end
		1'd1: begin
			sync_rhs_array_muxed10 <= videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			sync_rhs_array_muxed10 <= videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			sync_rhs_array_muxed10 <= videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed11 <= 1'd0;
	case (videosoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed11 <= videosoc_sdram_nop_we;
		end
		1'd1: begin
			sync_rhs_array_muxed11 <= videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			sync_rhs_array_muxed11 <= videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			sync_rhs_array_muxed11 <= videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed12 <= 1'd0;
	case (videosoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed12 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			sync_rhs_array_muxed12 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			sync_rhs_array_muxed12 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed13 <= 1'd0;
	case (videosoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed13 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed13 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			sync_rhs_array_muxed13 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			sync_rhs_array_muxed13 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed14 <= 15'd0;
	case (videosoc_sdram_sel2)
		1'd0: begin
			sync_rhs_array_muxed14 <= videosoc_sdram_nop_a;
		end
		1'd1: begin
			sync_rhs_array_muxed14 <= videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			sync_rhs_array_muxed14 <= videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			sync_rhs_array_muxed14 <= videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed15 <= 3'd0;
	case (videosoc_sdram_sel2)
		1'd0: begin
			sync_rhs_array_muxed15 <= videosoc_sdram_nop_ba;
		end
		1'd1: begin
			sync_rhs_array_muxed15 <= videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			sync_rhs_array_muxed15 <= videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			sync_rhs_array_muxed15 <= videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed16 <= 1'd0;
	case (videosoc_sdram_sel2)
		1'd0: begin
			sync_rhs_array_muxed16 <= videosoc_sdram_nop_cas;
		end
		1'd1: begin
			sync_rhs_array_muxed16 <= videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			sync_rhs_array_muxed16 <= videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			sync_rhs_array_muxed16 <= videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed17 <= 1'd0;
	case (videosoc_sdram_sel2)
		1'd0: begin
			sync_rhs_array_muxed17 <= videosoc_sdram_nop_ras;
		end
		1'd1: begin
			sync_rhs_array_muxed17 <= videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			sync_rhs_array_muxed17 <= videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			sync_rhs_array_muxed17 <= videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed18 <= 1'd0;
	case (videosoc_sdram_sel2)
		1'd0: begin
			sync_rhs_array_muxed18 <= videosoc_sdram_nop_we;
		end
		1'd1: begin
			sync_rhs_array_muxed18 <= videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			sync_rhs_array_muxed18 <= videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			sync_rhs_array_muxed18 <= videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed19 <= 1'd0;
	case (videosoc_sdram_sel2)
		1'd0: begin
			sync_rhs_array_muxed19 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed19 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			sync_rhs_array_muxed19 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			sync_rhs_array_muxed19 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed20 <= 1'd0;
	case (videosoc_sdram_sel2)
		1'd0: begin
			sync_rhs_array_muxed20 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed20 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			sync_rhs_array_muxed20 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			sync_rhs_array_muxed20 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed21 <= 15'd0;
	case (videosoc_sdram_sel3)
		1'd0: begin
			sync_rhs_array_muxed21 <= videosoc_sdram_nop_a;
		end
		1'd1: begin
			sync_rhs_array_muxed21 <= videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			sync_rhs_array_muxed21 <= videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			sync_rhs_array_muxed21 <= videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed22 <= 3'd0;
	case (videosoc_sdram_sel3)
		1'd0: begin
			sync_rhs_array_muxed22 <= videosoc_sdram_nop_ba;
		end
		1'd1: begin
			sync_rhs_array_muxed22 <= videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			sync_rhs_array_muxed22 <= videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			sync_rhs_array_muxed22 <= videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed23 <= 1'd0;
	case (videosoc_sdram_sel3)
		1'd0: begin
			sync_rhs_array_muxed23 <= videosoc_sdram_nop_cas;
		end
		1'd1: begin
			sync_rhs_array_muxed23 <= videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			sync_rhs_array_muxed23 <= videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			sync_rhs_array_muxed23 <= videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed24 <= 1'd0;
	case (videosoc_sdram_sel3)
		1'd0: begin
			sync_rhs_array_muxed24 <= videosoc_sdram_nop_ras;
		end
		1'd1: begin
			sync_rhs_array_muxed24 <= videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			sync_rhs_array_muxed24 <= videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			sync_rhs_array_muxed24 <= videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed25 <= 1'd0;
	case (videosoc_sdram_sel3)
		1'd0: begin
			sync_rhs_array_muxed25 <= videosoc_sdram_nop_we;
		end
		1'd1: begin
			sync_rhs_array_muxed25 <= videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			sync_rhs_array_muxed25 <= videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			sync_rhs_array_muxed25 <= videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed26 <= 1'd0;
	case (videosoc_sdram_sel3)
		1'd0: begin
			sync_rhs_array_muxed26 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed26 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			sync_rhs_array_muxed26 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			sync_rhs_array_muxed26 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	sync_rhs_array_muxed27 <= 1'd0;
	case (videosoc_sdram_sel3)
		1'd0: begin
			sync_rhs_array_muxed27 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed27 <= (videosoc_sdram_choose_cmd_cmd_valid & videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			sync_rhs_array_muxed27 <= (videosoc_sdram_choose_req_cmd_valid & videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			sync_rhs_array_muxed27 <= (videosoc_sdram_cmd_valid & videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
assign xilinxasyncresetsynchronizerimpl0 = ((~videosoc_pll_locked) | (~cpu_reset));
assign xilinxasyncresetsynchronizerimpl1 = ((~videosoc_pll_locked) | (~cpu_reset));
assign xilinxasyncresetsynchronizerimpl2 = ((~videosoc_pll_locked) | (~cpu_reset));
assign videosoc_uart_phy_rx = xilinxmultiregimpl0_regs1;
assign ethphy_status = xilinxmultiregimpl1_regs1;
assign ethmac_ps_preamble_error_toggle_o = xilinxmultiregimpl2_regs1;
assign ethmac_ps_crc_error_toggle_o = xilinxmultiregimpl3_regs1;
assign ethmac_tx_cdc_produce_rdomain = xilinxmultiregimpl4_regs1;
assign ethmac_tx_cdc_consume_wdomain = xilinxmultiregimpl5_regs1;
assign ethmac_rx_cdc_produce_rdomain = xilinxmultiregimpl6_regs1;
assign ethmac_rx_cdc_consume_wdomain = xilinxmultiregimpl7_regs1;
assign edid_scl_raw = xilinxmultiregimpl8_regs1;
assign edid_sda_raw = xilinxmultiregimpl9_regs1;
assign locked = xilinxmultiregimpl10_regs1;
assign xilinxasyncresetsynchronizerimpl5 = (~mmcm_locked);
assign xilinxasyncresetsynchronizerimpl6 = (~mmcm_locked);
assign s7datacapture0_do_delay_rst_toggle_o = xilinxmultiregimpl11_regs1;
assign s7datacapture0_do_delay_master_inc_toggle_o = xilinxmultiregimpl12_regs1;
assign s7datacapture0_do_delay_master_dec_toggle_o = xilinxmultiregimpl13_regs1;
assign s7datacapture0_do_delay_slave_inc_toggle_o = xilinxmultiregimpl14_regs1;
assign s7datacapture0_do_delay_slave_dec_toggle_o = xilinxmultiregimpl15_regs1;
assign s7datacapture0_status = xilinxmultiregimpl16_regs1;
assign s7datacapture0_do_reset_lateness_toggle_o = xilinxmultiregimpl17_regs1;
assign charsync0_char_synced_status = xilinxmultiregimpl18_regs1;
assign charsync0_ctl_pos_status = xilinxmultiregimpl19_regs1;
assign wer0_toggle_o = xilinxmultiregimpl20_regs1;
assign s7datacapture1_do_delay_rst_toggle_o = xilinxmultiregimpl21_regs1;
assign s7datacapture1_do_delay_master_inc_toggle_o = xilinxmultiregimpl22_regs1;
assign s7datacapture1_do_delay_master_dec_toggle_o = xilinxmultiregimpl23_regs1;
assign s7datacapture1_do_delay_slave_inc_toggle_o = xilinxmultiregimpl24_regs1;
assign s7datacapture1_do_delay_slave_dec_toggle_o = xilinxmultiregimpl25_regs1;
assign s7datacapture1_status = xilinxmultiregimpl26_regs1;
assign s7datacapture1_do_reset_lateness_toggle_o = xilinxmultiregimpl27_regs1;
assign charsync1_char_synced_status = xilinxmultiregimpl28_regs1;
assign charsync1_ctl_pos_status = xilinxmultiregimpl29_regs1;
assign wer1_toggle_o = xilinxmultiregimpl30_regs1;
assign s7datacapture2_do_delay_rst_toggle_o = xilinxmultiregimpl31_regs1;
assign s7datacapture2_do_delay_master_inc_toggle_o = xilinxmultiregimpl32_regs1;
assign s7datacapture2_do_delay_master_dec_toggle_o = xilinxmultiregimpl33_regs1;
assign s7datacapture2_do_delay_slave_inc_toggle_o = xilinxmultiregimpl34_regs1;
assign s7datacapture2_do_delay_slave_dec_toggle_o = xilinxmultiregimpl35_regs1;
assign s7datacapture2_status = xilinxmultiregimpl36_regs1;
assign s7datacapture2_do_reset_lateness_toggle_o = xilinxmultiregimpl37_regs1;
assign charsync2_char_synced_status = xilinxmultiregimpl38_regs1;
assign charsync2_ctl_pos_status = xilinxmultiregimpl39_regs1;
assign wer2_toggle_o = xilinxmultiregimpl40_regs1;
assign chansync_status = xilinxmultiregimpl41_regs1;
assign resdetection_hres_status = xilinxmultiregimpl42_regs1;
assign resdetection_vres_status = xilinxmultiregimpl43_regs1;
assign frame_fifo_produce_rdomain = xilinxmultiregimpl44_regs1;
assign frame_fifo_consume_wdomain = xilinxmultiregimpl45_regs1;
assign frame_sys_overflow = xilinxmultiregimpl46_regs1;
assign frame_overflow_reset_toggle_o = xilinxmultiregimpl47_regs1;
assign frame_overflow_reset_ack_toggle_o = xilinxmultiregimpl48_regs1;
assign hdmi_in0_freq_gray_decoder_i = xilinxmultiregimpl49_regs1;
assign hdmi_out0_dram_port_cmd_fifo_produce_rdomain = xilinxmultiregimpl50_regs1;
assign hdmi_out0_dram_port_cmd_fifo_consume_wdomain = xilinxmultiregimpl51_regs1;
assign hdmi_out0_dram_port_rdata_fifo_produce_rdomain = xilinxmultiregimpl52_regs1;
assign hdmi_out0_dram_port_rdata_fifo_consume_wdomain = xilinxmultiregimpl53_regs1;
assign hdmi_out0_core_initiator_cdc_produce_rdomain = xilinxmultiregimpl54_regs1;
assign hdmi_out0_core_initiator_cdc_consume_wdomain = xilinxmultiregimpl55_regs1;
assign hdmi_out0_core_underflow_enable = xilinxmultiregimpl56_regs1;
assign hdmi_out0_core_toggle_o = xilinxmultiregimpl57_regs1;

always @(posedge clk200_clk) begin
	if ((videosoc_reset_counter != 1'd0)) begin
		videosoc_reset_counter <= (videosoc_reset_counter - 1'd1);
	end else begin
		videosoc_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		videosoc_reset_counter <= 4'd15;
		videosoc_ic_reset <= 1'd1;
	end
end

always @(posedge data0_cap_read_clk) begin
	if ((s7datacapture0_gearbox_rdpointer == 3'd7)) begin
		s7datacapture0_gearbox_rdpointer <= 1'd0;
	end else begin
		s7datacapture0_gearbox_rdpointer <= (s7datacapture0_gearbox_rdpointer + 1'd1);
	end
	case (s7datacapture0_gearbox_rdpointer)
		1'd0: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[9:0];
		end
		1'd1: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[19:10];
		end
		2'd2: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[29:20];
		end
		2'd3: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[39:30];
		end
		3'd4: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[49:40];
		end
		3'd5: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[59:50];
		end
		3'd6: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[69:60];
		end
		3'd7: begin
			s7datacapture0_gearbox_o <= s7datacapture0_gearbox_storage[79:70];
		end
	endcase
	if (data0_cap_read_rst) begin
		s7datacapture0_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge data0_cap_write_clk) begin
	if ((s7datacapture0_gearbox_wrpointer == 4'd9)) begin
		s7datacapture0_gearbox_wrpointer <= 1'd0;
	end else begin
		s7datacapture0_gearbox_wrpointer <= (s7datacapture0_gearbox_wrpointer + 1'd1);
	end
	case (s7datacapture0_gearbox_wrpointer)
		1'd0: begin
			s7datacapture0_gearbox_storage[7:0] <= s7datacapture0_gearbox_i;
		end
		1'd1: begin
			s7datacapture0_gearbox_storage[15:8] <= s7datacapture0_gearbox_i;
		end
		2'd2: begin
			s7datacapture0_gearbox_storage[23:16] <= s7datacapture0_gearbox_i;
		end
		2'd3: begin
			s7datacapture0_gearbox_storage[31:24] <= s7datacapture0_gearbox_i;
		end
		3'd4: begin
			s7datacapture0_gearbox_storage[39:32] <= s7datacapture0_gearbox_i;
		end
		3'd5: begin
			s7datacapture0_gearbox_storage[47:40] <= s7datacapture0_gearbox_i;
		end
		3'd6: begin
			s7datacapture0_gearbox_storage[55:48] <= s7datacapture0_gearbox_i;
		end
		3'd7: begin
			s7datacapture0_gearbox_storage[63:56] <= s7datacapture0_gearbox_i;
		end
		4'd8: begin
			s7datacapture0_gearbox_storage[71:64] <= s7datacapture0_gearbox_i;
		end
		4'd9: begin
			s7datacapture0_gearbox_storage[79:72] <= s7datacapture0_gearbox_i;
		end
	endcase
	if (data0_cap_write_rst) begin
		s7datacapture0_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge data1_cap_read_clk) begin
	if ((s7datacapture1_gearbox_rdpointer == 3'd7)) begin
		s7datacapture1_gearbox_rdpointer <= 1'd0;
	end else begin
		s7datacapture1_gearbox_rdpointer <= (s7datacapture1_gearbox_rdpointer + 1'd1);
	end
	case (s7datacapture1_gearbox_rdpointer)
		1'd0: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[9:0];
		end
		1'd1: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[19:10];
		end
		2'd2: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[29:20];
		end
		2'd3: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[39:30];
		end
		3'd4: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[49:40];
		end
		3'd5: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[59:50];
		end
		3'd6: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[69:60];
		end
		3'd7: begin
			s7datacapture1_gearbox_o <= s7datacapture1_gearbox_storage[79:70];
		end
	endcase
	if (data1_cap_read_rst) begin
		s7datacapture1_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge data1_cap_write_clk) begin
	if ((s7datacapture1_gearbox_wrpointer == 4'd9)) begin
		s7datacapture1_gearbox_wrpointer <= 1'd0;
	end else begin
		s7datacapture1_gearbox_wrpointer <= (s7datacapture1_gearbox_wrpointer + 1'd1);
	end
	case (s7datacapture1_gearbox_wrpointer)
		1'd0: begin
			s7datacapture1_gearbox_storage[7:0] <= s7datacapture1_gearbox_i;
		end
		1'd1: begin
			s7datacapture1_gearbox_storage[15:8] <= s7datacapture1_gearbox_i;
		end
		2'd2: begin
			s7datacapture1_gearbox_storage[23:16] <= s7datacapture1_gearbox_i;
		end
		2'd3: begin
			s7datacapture1_gearbox_storage[31:24] <= s7datacapture1_gearbox_i;
		end
		3'd4: begin
			s7datacapture1_gearbox_storage[39:32] <= s7datacapture1_gearbox_i;
		end
		3'd5: begin
			s7datacapture1_gearbox_storage[47:40] <= s7datacapture1_gearbox_i;
		end
		3'd6: begin
			s7datacapture1_gearbox_storage[55:48] <= s7datacapture1_gearbox_i;
		end
		3'd7: begin
			s7datacapture1_gearbox_storage[63:56] <= s7datacapture1_gearbox_i;
		end
		4'd8: begin
			s7datacapture1_gearbox_storage[71:64] <= s7datacapture1_gearbox_i;
		end
		4'd9: begin
			s7datacapture1_gearbox_storage[79:72] <= s7datacapture1_gearbox_i;
		end
	endcase
	if (data1_cap_write_rst) begin
		s7datacapture1_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge data2_cap_read_clk) begin
	if ((s7datacapture2_gearbox_rdpointer == 3'd7)) begin
		s7datacapture2_gearbox_rdpointer <= 1'd0;
	end else begin
		s7datacapture2_gearbox_rdpointer <= (s7datacapture2_gearbox_rdpointer + 1'd1);
	end
	case (s7datacapture2_gearbox_rdpointer)
		1'd0: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[9:0];
		end
		1'd1: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[19:10];
		end
		2'd2: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[29:20];
		end
		2'd3: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[39:30];
		end
		3'd4: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[49:40];
		end
		3'd5: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[59:50];
		end
		3'd6: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[69:60];
		end
		3'd7: begin
			s7datacapture2_gearbox_o <= s7datacapture2_gearbox_storage[79:70];
		end
	endcase
	if (data2_cap_read_rst) begin
		s7datacapture2_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge data2_cap_write_clk) begin
	if ((s7datacapture2_gearbox_wrpointer == 4'd9)) begin
		s7datacapture2_gearbox_wrpointer <= 1'd0;
	end else begin
		s7datacapture2_gearbox_wrpointer <= (s7datacapture2_gearbox_wrpointer + 1'd1);
	end
	case (s7datacapture2_gearbox_wrpointer)
		1'd0: begin
			s7datacapture2_gearbox_storage[7:0] <= s7datacapture2_gearbox_i;
		end
		1'd1: begin
			s7datacapture2_gearbox_storage[15:8] <= s7datacapture2_gearbox_i;
		end
		2'd2: begin
			s7datacapture2_gearbox_storage[23:16] <= s7datacapture2_gearbox_i;
		end
		2'd3: begin
			s7datacapture2_gearbox_storage[31:24] <= s7datacapture2_gearbox_i;
		end
		3'd4: begin
			s7datacapture2_gearbox_storage[39:32] <= s7datacapture2_gearbox_i;
		end
		3'd5: begin
			s7datacapture2_gearbox_storage[47:40] <= s7datacapture2_gearbox_i;
		end
		3'd6: begin
			s7datacapture2_gearbox_storage[55:48] <= s7datacapture2_gearbox_i;
		end
		3'd7: begin
			s7datacapture2_gearbox_storage[63:56] <= s7datacapture2_gearbox_i;
		end
		4'd8: begin
			s7datacapture2_gearbox_storage[71:64] <= s7datacapture2_gearbox_i;
		end
		4'd9: begin
			s7datacapture2_gearbox_storage[79:72] <= s7datacapture2_gearbox_i;
		end
	endcase
	if (data2_cap_write_rst) begin
		s7datacapture2_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge eth_rx_clk) begin
	ethphy_rx_ctl_d <= ethphy_rx_ctl;
	ethphy_source_valid <= ethphy_rx_ctl;
	ethphy_source_payload_data <= ethphy_rx_data;
	liteethmacpreamblechecker_state <= liteethmacpreamblechecker_next_state;
	if (ethmac_crc32_checker_crc_ce) begin
		ethmac_crc32_checker_crc_reg <= ethmac_crc32_checker_crc_next;
	end
	if (ethmac_crc32_checker_crc_reset) begin
		ethmac_crc32_checker_crc_reg <= 32'd4294967295;
	end
	if (((ethmac_crc32_checker_syncfifo_syncfifo_we & ethmac_crc32_checker_syncfifo_syncfifo_writable) & (~ethmac_crc32_checker_syncfifo_replace))) begin
		if ((ethmac_crc32_checker_syncfifo_produce == 3'd4)) begin
			ethmac_crc32_checker_syncfifo_produce <= 1'd0;
		end else begin
			ethmac_crc32_checker_syncfifo_produce <= (ethmac_crc32_checker_syncfifo_produce + 1'd1);
		end
	end
	if (ethmac_crc32_checker_syncfifo_do_read) begin
		if ((ethmac_crc32_checker_syncfifo_consume == 3'd4)) begin
			ethmac_crc32_checker_syncfifo_consume <= 1'd0;
		end else begin
			ethmac_crc32_checker_syncfifo_consume <= (ethmac_crc32_checker_syncfifo_consume + 1'd1);
		end
	end
	if (((ethmac_crc32_checker_syncfifo_syncfifo_we & ethmac_crc32_checker_syncfifo_syncfifo_writable) & (~ethmac_crc32_checker_syncfifo_replace))) begin
		if ((~ethmac_crc32_checker_syncfifo_do_read)) begin
			ethmac_crc32_checker_syncfifo_level <= (ethmac_crc32_checker_syncfifo_level + 1'd1);
		end
	end else begin
		if (ethmac_crc32_checker_syncfifo_do_read) begin
			ethmac_crc32_checker_syncfifo_level <= (ethmac_crc32_checker_syncfifo_level - 1'd1);
		end
	end
	if (ethmac_crc32_checker_fifo_reset) begin
		ethmac_crc32_checker_syncfifo_level <= 3'd0;
		ethmac_crc32_checker_syncfifo_produce <= 3'd0;
		ethmac_crc32_checker_syncfifo_consume <= 3'd0;
	end
	liteethmaccrc32checker_state <= liteethmaccrc32checker_next_state;
	if (ethmac_ps_preamble_error_i) begin
		ethmac_ps_preamble_error_toggle_i <= (~ethmac_ps_preamble_error_toggle_i);
	end
	if (ethmac_ps_crc_error_i) begin
		ethmac_ps_crc_error_toggle_i <= (~ethmac_ps_crc_error_toggle_i);
	end
	if (ethmac_rx_converter_converter_source_ready) begin
		ethmac_rx_converter_converter_strobe_all <= 1'd0;
	end
	if (ethmac_rx_converter_converter_load_part) begin
		if (((ethmac_rx_converter_converter_demux == 2'd3) | ethmac_rx_converter_converter_sink_last)) begin
			ethmac_rx_converter_converter_demux <= 1'd0;
			ethmac_rx_converter_converter_strobe_all <= 1'd1;
		end else begin
			ethmac_rx_converter_converter_demux <= (ethmac_rx_converter_converter_demux + 1'd1);
		end
	end
	if ((ethmac_rx_converter_converter_source_valid & ethmac_rx_converter_converter_source_ready)) begin
		if ((ethmac_rx_converter_converter_sink_valid & ethmac_rx_converter_converter_sink_ready)) begin
			ethmac_rx_converter_converter_source_first <= ethmac_rx_converter_converter_sink_first;
			ethmac_rx_converter_converter_source_last <= ethmac_rx_converter_converter_sink_last;
		end else begin
			ethmac_rx_converter_converter_source_first <= 1'd0;
			ethmac_rx_converter_converter_source_last <= 1'd0;
		end
	end else begin
		if ((ethmac_rx_converter_converter_sink_valid & ethmac_rx_converter_converter_sink_ready)) begin
			ethmac_rx_converter_converter_source_first <= (ethmac_rx_converter_converter_sink_first | ethmac_rx_converter_converter_source_first);
			ethmac_rx_converter_converter_source_last <= (ethmac_rx_converter_converter_sink_last | ethmac_rx_converter_converter_source_last);
		end
	end
	if (ethmac_rx_converter_converter_load_part) begin
		case (ethmac_rx_converter_converter_demux)
			1'd0: begin
				ethmac_rx_converter_converter_source_payload_data[39:30] <= ethmac_rx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				ethmac_rx_converter_converter_source_payload_data[29:20] <= ethmac_rx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				ethmac_rx_converter_converter_source_payload_data[19:10] <= ethmac_rx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				ethmac_rx_converter_converter_source_payload_data[9:0] <= ethmac_rx_converter_converter_sink_payload_data;
			end
		endcase
	end
	if (ethmac_rx_converter_converter_load_part) begin
		ethmac_rx_converter_converter_source_payload_valid_token_count <= (ethmac_rx_converter_converter_demux + 1'd1);
	end
	ethmac_rx_cdc_graycounter0_q_binary <= ethmac_rx_cdc_graycounter0_q_next_binary;
	ethmac_rx_cdc_graycounter0_q <= ethmac_rx_cdc_graycounter0_q_next;
	if (eth_rx_rst) begin
		ethphy_source_valid <= 1'd0;
		ethphy_rx_ctl_d <= 1'd0;
		ethmac_crc32_checker_crc_reg <= 32'd4294967295;
		ethmac_crc32_checker_syncfifo_level <= 3'd0;
		ethmac_crc32_checker_syncfifo_produce <= 3'd0;
		ethmac_crc32_checker_syncfifo_consume <= 3'd0;
		ethmac_rx_converter_converter_source_first <= 1'd0;
		ethmac_rx_converter_converter_source_last <= 1'd0;
		ethmac_rx_converter_converter_demux <= 2'd0;
		ethmac_rx_converter_converter_strobe_all <= 1'd0;
		ethmac_rx_cdc_graycounter0_q <= 7'd0;
		ethmac_rx_cdc_graycounter0_q_binary <= 7'd0;
		liteethmacpreamblechecker_state <= 1'd0;
		liteethmaccrc32checker_state <= 2'd0;
	end
	xilinxmultiregimpl7_regs0 <= ethmac_rx_cdc_graycounter1_q;
	xilinxmultiregimpl7_regs1 <= xilinxmultiregimpl7_regs0;
end

always @(posedge eth_tx_clk) begin
	if (ethmac_tx_gap_inserter_counter_reset) begin
		ethmac_tx_gap_inserter_counter <= 1'd0;
	end else begin
		if (ethmac_tx_gap_inserter_counter_ce) begin
			ethmac_tx_gap_inserter_counter <= (ethmac_tx_gap_inserter_counter + 1'd1);
		end
	end
	liteethmacgap_state <= liteethmacgap_next_state;
	if (ethmac_preamble_inserter_clr_cnt) begin
		ethmac_preamble_inserter_cnt <= 1'd0;
	end else begin
		if (ethmac_preamble_inserter_inc_cnt) begin
			ethmac_preamble_inserter_cnt <= (ethmac_preamble_inserter_cnt + 1'd1);
		end
	end
	liteethmacpreambleinserter_state <= liteethmacpreambleinserter_next_state;
	if (ethmac_crc32_inserter_is_ongoing0) begin
		ethmac_crc32_inserter_cnt <= 2'd3;
	end else begin
		if ((ethmac_crc32_inserter_is_ongoing1 & (~ethmac_crc32_inserter_cnt_done))) begin
			ethmac_crc32_inserter_cnt <= (ethmac_crc32_inserter_cnt - ethmac_crc32_inserter_source_ready);
		end
	end
	if (ethmac_crc32_inserter_ce) begin
		ethmac_crc32_inserter_reg <= ethmac_crc32_inserter_next;
	end
	if (ethmac_crc32_inserter_reset) begin
		ethmac_crc32_inserter_reg <= 32'd4294967295;
	end
	liteethmaccrc32inserter_state <= liteethmaccrc32inserter_next_state;
	if (ethmac_padding_inserter_counter_reset) begin
		ethmac_padding_inserter_counter <= 1'd0;
	end else begin
		if (ethmac_padding_inserter_counter_ce) begin
			ethmac_padding_inserter_counter <= (ethmac_padding_inserter_counter + 1'd1);
		end
	end
	liteethmacpaddinginserter_state <= liteethmacpaddinginserter_next_state;
	if ((ethmac_tx_last_be_sink_valid & ethmac_tx_last_be_sink_ready)) begin
		if (ethmac_tx_last_be_sink_last) begin
			ethmac_tx_last_be_ongoing <= 1'd1;
		end else begin
			if (ethmac_tx_last_be_sink_payload_last_be) begin
				ethmac_tx_last_be_ongoing <= 1'd0;
			end
		end
	end
	if ((ethmac_tx_converter_converter_source_valid & ethmac_tx_converter_converter_source_ready)) begin
		if (ethmac_tx_converter_converter_last) begin
			ethmac_tx_converter_converter_mux <= 1'd0;
		end else begin
			ethmac_tx_converter_converter_mux <= (ethmac_tx_converter_converter_mux + 1'd1);
		end
	end
	ethmac_tx_cdc_graycounter1_q_binary <= ethmac_tx_cdc_graycounter1_q_next_binary;
	ethmac_tx_cdc_graycounter1_q <= ethmac_tx_cdc_graycounter1_q_next;
	if (eth_tx_rst) begin
		ethmac_crc32_inserter_reg <= 32'd4294967295;
		ethmac_crc32_inserter_cnt <= 2'd3;
		ethmac_padding_inserter_counter <= 16'd1;
		ethmac_tx_last_be_ongoing <= 1'd1;
		ethmac_tx_converter_converter_mux <= 2'd0;
		ethmac_tx_cdc_graycounter1_q <= 7'd0;
		ethmac_tx_cdc_graycounter1_q_binary <= 7'd0;
		liteethmacgap_state <= 1'd0;
		liteethmacpreambleinserter_state <= 2'd0;
		liteethmaccrc32inserter_state <= 2'd0;
		liteethmacpaddinginserter_state <= 1'd0;
	end
	xilinxmultiregimpl4_regs0 <= ethmac_tx_cdc_graycounter0_q;
	xilinxmultiregimpl4_regs1 <= xilinxmultiregimpl4_regs0;
end

always @(posedge fmeter_clk) begin
	hdmi_in0_freq_q_binary <= hdmi_in0_freq_q_next_binary;
	hdmi_in0_freq_q <= hdmi_in0_freq_q_next;
end

always @(posedge hdmi_in0_pix_clk) begin
	charsync0_raw_data1 <= charsync0_raw_data;
	charsync0_found_control <= 1'd0;
	if (((((charsync0_raw[9:0] == 10'd852) | (charsync0_raw[9:0] == 8'd171)) | (charsync0_raw[9:0] == 9'd340)) | (charsync0_raw[9:0] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 1'd0;
	end
	if (((((charsync0_raw[10:1] == 10'd852) | (charsync0_raw[10:1] == 8'd171)) | (charsync0_raw[10:1] == 9'd340)) | (charsync0_raw[10:1] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 1'd1;
	end
	if (((((charsync0_raw[11:2] == 10'd852) | (charsync0_raw[11:2] == 8'd171)) | (charsync0_raw[11:2] == 9'd340)) | (charsync0_raw[11:2] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 2'd2;
	end
	if (((((charsync0_raw[12:3] == 10'd852) | (charsync0_raw[12:3] == 8'd171)) | (charsync0_raw[12:3] == 9'd340)) | (charsync0_raw[12:3] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 2'd3;
	end
	if (((((charsync0_raw[13:4] == 10'd852) | (charsync0_raw[13:4] == 8'd171)) | (charsync0_raw[13:4] == 9'd340)) | (charsync0_raw[13:4] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 3'd4;
	end
	if (((((charsync0_raw[14:5] == 10'd852) | (charsync0_raw[14:5] == 8'd171)) | (charsync0_raw[14:5] == 9'd340)) | (charsync0_raw[14:5] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 3'd5;
	end
	if (((((charsync0_raw[15:6] == 10'd852) | (charsync0_raw[15:6] == 8'd171)) | (charsync0_raw[15:6] == 9'd340)) | (charsync0_raw[15:6] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 3'd6;
	end
	if (((((charsync0_raw[16:7] == 10'd852) | (charsync0_raw[16:7] == 8'd171)) | (charsync0_raw[16:7] == 9'd340)) | (charsync0_raw[16:7] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 3'd7;
	end
	if (((((charsync0_raw[17:8] == 10'd852) | (charsync0_raw[17:8] == 8'd171)) | (charsync0_raw[17:8] == 9'd340)) | (charsync0_raw[17:8] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 4'd8;
	end
	if (((((charsync0_raw[18:9] == 10'd852) | (charsync0_raw[18:9] == 8'd171)) | (charsync0_raw[18:9] == 9'd340)) | (charsync0_raw[18:9] == 10'd683))) begin
		charsync0_found_control <= 1'd1;
		charsync0_control_position <= 4'd9;
	end
	if ((charsync0_found_control & (charsync0_control_position == charsync0_previous_control_position))) begin
		if ((charsync0_control_counter == 3'd7)) begin
			charsync0_control_counter <= 1'd0;
			charsync0_synced <= 1'd1;
			charsync0_word_sel <= charsync0_control_position;
		end else begin
			charsync0_control_counter <= (charsync0_control_counter + 1'd1);
		end
	end else begin
		charsync0_control_counter <= 1'd0;
	end
	charsync0_previous_control_position <= charsync0_control_position;
	charsync0_data <= (charsync0_raw >>> charsync0_word_sel);
	wer0_data_r <= wer0_data[8:0];
	wer0_transition_count <= (((((((wer0_transitions[0] + wer0_transitions[1]) + wer0_transitions[2]) + wer0_transitions[3]) + wer0_transitions[4]) + wer0_transitions[5]) + wer0_transitions[6]) + wer0_transitions[7]);
	wer0_is_control <= ((((wer0_data_r == 10'd852) | (wer0_data_r == 8'd171)) | (wer0_data_r == 9'd340)) | (wer0_data_r == 10'd683));
	wer0_is_error <= ((wer0_transition_count > 3'd4) & (~wer0_is_control));
	{wer0_period_done, wer0_period_counter} <= (wer0_period_counter + 1'd1);
	wer0_wer_counter_r_updated <= wer0_period_done;
	if (wer0_period_done) begin
		wer0_wer_counter_r <= wer0_wer_counter;
		wer0_wer_counter <= 1'd0;
	end else begin
		if (wer0_is_error) begin
			wer0_wer_counter <= (wer0_wer_counter + 1'd1);
		end
	end
	if (wer0_i) begin
		wer0_toggle_i <= (~wer0_toggle_i);
	end
	decoding0_output_de <= 1'd1;
	if ((decoding0_input == 10'd852)) begin
		decoding0_output_de <= 1'd0;
		decoding0_output_c <= 1'd0;
	end
	if ((decoding0_input == 8'd171)) begin
		decoding0_output_de <= 1'd0;
		decoding0_output_c <= 1'd1;
	end
	if ((decoding0_input == 9'd340)) begin
		decoding0_output_de <= 1'd0;
		decoding0_output_c <= 2'd2;
	end
	if ((decoding0_input == 10'd683)) begin
		decoding0_output_de <= 1'd0;
		decoding0_output_c <= 2'd3;
	end
	decoding0_output_d[0] <= (decoding0_input[0] ^ decoding0_input[9]);
	decoding0_output_d[1] <= ((decoding0_input[1] ^ decoding0_input[0]) ^ (~decoding0_input[8]));
	decoding0_output_d[2] <= ((decoding0_input[2] ^ decoding0_input[1]) ^ (~decoding0_input[8]));
	decoding0_output_d[3] <= ((decoding0_input[3] ^ decoding0_input[2]) ^ (~decoding0_input[8]));
	decoding0_output_d[4] <= ((decoding0_input[4] ^ decoding0_input[3]) ^ (~decoding0_input[8]));
	decoding0_output_d[5] <= ((decoding0_input[5] ^ decoding0_input[4]) ^ (~decoding0_input[8]));
	decoding0_output_d[6] <= ((decoding0_input[6] ^ decoding0_input[5]) ^ (~decoding0_input[8]));
	decoding0_output_d[7] <= ((decoding0_input[7] ^ decoding0_input[6]) ^ (~decoding0_input[8]));
	decoding0_valid_o <= decoding0_valid_i;
	charsync1_raw_data1 <= charsync1_raw_data;
	charsync1_found_control <= 1'd0;
	if (((((charsync1_raw[9:0] == 10'd852) | (charsync1_raw[9:0] == 8'd171)) | (charsync1_raw[9:0] == 9'd340)) | (charsync1_raw[9:0] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 1'd0;
	end
	if (((((charsync1_raw[10:1] == 10'd852) | (charsync1_raw[10:1] == 8'd171)) | (charsync1_raw[10:1] == 9'd340)) | (charsync1_raw[10:1] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 1'd1;
	end
	if (((((charsync1_raw[11:2] == 10'd852) | (charsync1_raw[11:2] == 8'd171)) | (charsync1_raw[11:2] == 9'd340)) | (charsync1_raw[11:2] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 2'd2;
	end
	if (((((charsync1_raw[12:3] == 10'd852) | (charsync1_raw[12:3] == 8'd171)) | (charsync1_raw[12:3] == 9'd340)) | (charsync1_raw[12:3] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 2'd3;
	end
	if (((((charsync1_raw[13:4] == 10'd852) | (charsync1_raw[13:4] == 8'd171)) | (charsync1_raw[13:4] == 9'd340)) | (charsync1_raw[13:4] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 3'd4;
	end
	if (((((charsync1_raw[14:5] == 10'd852) | (charsync1_raw[14:5] == 8'd171)) | (charsync1_raw[14:5] == 9'd340)) | (charsync1_raw[14:5] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 3'd5;
	end
	if (((((charsync1_raw[15:6] == 10'd852) | (charsync1_raw[15:6] == 8'd171)) | (charsync1_raw[15:6] == 9'd340)) | (charsync1_raw[15:6] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 3'd6;
	end
	if (((((charsync1_raw[16:7] == 10'd852) | (charsync1_raw[16:7] == 8'd171)) | (charsync1_raw[16:7] == 9'd340)) | (charsync1_raw[16:7] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 3'd7;
	end
	if (((((charsync1_raw[17:8] == 10'd852) | (charsync1_raw[17:8] == 8'd171)) | (charsync1_raw[17:8] == 9'd340)) | (charsync1_raw[17:8] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 4'd8;
	end
	if (((((charsync1_raw[18:9] == 10'd852) | (charsync1_raw[18:9] == 8'd171)) | (charsync1_raw[18:9] == 9'd340)) | (charsync1_raw[18:9] == 10'd683))) begin
		charsync1_found_control <= 1'd1;
		charsync1_control_position <= 4'd9;
	end
	if ((charsync1_found_control & (charsync1_control_position == charsync1_previous_control_position))) begin
		if ((charsync1_control_counter == 3'd7)) begin
			charsync1_control_counter <= 1'd0;
			charsync1_synced <= 1'd1;
			charsync1_word_sel <= charsync1_control_position;
		end else begin
			charsync1_control_counter <= (charsync1_control_counter + 1'd1);
		end
	end else begin
		charsync1_control_counter <= 1'd0;
	end
	charsync1_previous_control_position <= charsync1_control_position;
	charsync1_data <= (charsync1_raw >>> charsync1_word_sel);
	wer1_data_r <= wer1_data[8:0];
	wer1_transition_count <= (((((((wer1_transitions[0] + wer1_transitions[1]) + wer1_transitions[2]) + wer1_transitions[3]) + wer1_transitions[4]) + wer1_transitions[5]) + wer1_transitions[6]) + wer1_transitions[7]);
	wer1_is_control <= ((((wer1_data_r == 10'd852) | (wer1_data_r == 8'd171)) | (wer1_data_r == 9'd340)) | (wer1_data_r == 10'd683));
	wer1_is_error <= ((wer1_transition_count > 3'd4) & (~wer1_is_control));
	{wer1_period_done, wer1_period_counter} <= (wer1_period_counter + 1'd1);
	wer1_wer_counter_r_updated <= wer1_period_done;
	if (wer1_period_done) begin
		wer1_wer_counter_r <= wer1_wer_counter;
		wer1_wer_counter <= 1'd0;
	end else begin
		if (wer1_is_error) begin
			wer1_wer_counter <= (wer1_wer_counter + 1'd1);
		end
	end
	if (wer1_i) begin
		wer1_toggle_i <= (~wer1_toggle_i);
	end
	decoding1_output_de <= 1'd1;
	if ((decoding1_input == 10'd852)) begin
		decoding1_output_de <= 1'd0;
		decoding1_output_c <= 1'd0;
	end
	if ((decoding1_input == 8'd171)) begin
		decoding1_output_de <= 1'd0;
		decoding1_output_c <= 1'd1;
	end
	if ((decoding1_input == 9'd340)) begin
		decoding1_output_de <= 1'd0;
		decoding1_output_c <= 2'd2;
	end
	if ((decoding1_input == 10'd683)) begin
		decoding1_output_de <= 1'd0;
		decoding1_output_c <= 2'd3;
	end
	decoding1_output_d[0] <= (decoding1_input[0] ^ decoding1_input[9]);
	decoding1_output_d[1] <= ((decoding1_input[1] ^ decoding1_input[0]) ^ (~decoding1_input[8]));
	decoding1_output_d[2] <= ((decoding1_input[2] ^ decoding1_input[1]) ^ (~decoding1_input[8]));
	decoding1_output_d[3] <= ((decoding1_input[3] ^ decoding1_input[2]) ^ (~decoding1_input[8]));
	decoding1_output_d[4] <= ((decoding1_input[4] ^ decoding1_input[3]) ^ (~decoding1_input[8]));
	decoding1_output_d[5] <= ((decoding1_input[5] ^ decoding1_input[4]) ^ (~decoding1_input[8]));
	decoding1_output_d[6] <= ((decoding1_input[6] ^ decoding1_input[5]) ^ (~decoding1_input[8]));
	decoding1_output_d[7] <= ((decoding1_input[7] ^ decoding1_input[6]) ^ (~decoding1_input[8]));
	decoding1_valid_o <= decoding1_valid_i;
	charsync2_raw_data1 <= charsync2_raw_data;
	charsync2_found_control <= 1'd0;
	if (((((charsync2_raw[9:0] == 10'd852) | (charsync2_raw[9:0] == 8'd171)) | (charsync2_raw[9:0] == 9'd340)) | (charsync2_raw[9:0] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 1'd0;
	end
	if (((((charsync2_raw[10:1] == 10'd852) | (charsync2_raw[10:1] == 8'd171)) | (charsync2_raw[10:1] == 9'd340)) | (charsync2_raw[10:1] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 1'd1;
	end
	if (((((charsync2_raw[11:2] == 10'd852) | (charsync2_raw[11:2] == 8'd171)) | (charsync2_raw[11:2] == 9'd340)) | (charsync2_raw[11:2] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 2'd2;
	end
	if (((((charsync2_raw[12:3] == 10'd852) | (charsync2_raw[12:3] == 8'd171)) | (charsync2_raw[12:3] == 9'd340)) | (charsync2_raw[12:3] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 2'd3;
	end
	if (((((charsync2_raw[13:4] == 10'd852) | (charsync2_raw[13:4] == 8'd171)) | (charsync2_raw[13:4] == 9'd340)) | (charsync2_raw[13:4] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 3'd4;
	end
	if (((((charsync2_raw[14:5] == 10'd852) | (charsync2_raw[14:5] == 8'd171)) | (charsync2_raw[14:5] == 9'd340)) | (charsync2_raw[14:5] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 3'd5;
	end
	if (((((charsync2_raw[15:6] == 10'd852) | (charsync2_raw[15:6] == 8'd171)) | (charsync2_raw[15:6] == 9'd340)) | (charsync2_raw[15:6] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 3'd6;
	end
	if (((((charsync2_raw[16:7] == 10'd852) | (charsync2_raw[16:7] == 8'd171)) | (charsync2_raw[16:7] == 9'd340)) | (charsync2_raw[16:7] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 3'd7;
	end
	if (((((charsync2_raw[17:8] == 10'd852) | (charsync2_raw[17:8] == 8'd171)) | (charsync2_raw[17:8] == 9'd340)) | (charsync2_raw[17:8] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 4'd8;
	end
	if (((((charsync2_raw[18:9] == 10'd852) | (charsync2_raw[18:9] == 8'd171)) | (charsync2_raw[18:9] == 9'd340)) | (charsync2_raw[18:9] == 10'd683))) begin
		charsync2_found_control <= 1'd1;
		charsync2_control_position <= 4'd9;
	end
	if ((charsync2_found_control & (charsync2_control_position == charsync2_previous_control_position))) begin
		if ((charsync2_control_counter == 3'd7)) begin
			charsync2_control_counter <= 1'd0;
			charsync2_synced <= 1'd1;
			charsync2_word_sel <= charsync2_control_position;
		end else begin
			charsync2_control_counter <= (charsync2_control_counter + 1'd1);
		end
	end else begin
		charsync2_control_counter <= 1'd0;
	end
	charsync2_previous_control_position <= charsync2_control_position;
	charsync2_data <= (charsync2_raw >>> charsync2_word_sel);
	wer2_data_r <= wer2_data[8:0];
	wer2_transition_count <= (((((((wer2_transitions[0] + wer2_transitions[1]) + wer2_transitions[2]) + wer2_transitions[3]) + wer2_transitions[4]) + wer2_transitions[5]) + wer2_transitions[6]) + wer2_transitions[7]);
	wer2_is_control <= ((((wer2_data_r == 10'd852) | (wer2_data_r == 8'd171)) | (wer2_data_r == 9'd340)) | (wer2_data_r == 10'd683));
	wer2_is_error <= ((wer2_transition_count > 3'd4) & (~wer2_is_control));
	{wer2_period_done, wer2_period_counter} <= (wer2_period_counter + 1'd1);
	wer2_wer_counter_r_updated <= wer2_period_done;
	if (wer2_period_done) begin
		wer2_wer_counter_r <= wer2_wer_counter;
		wer2_wer_counter <= 1'd0;
	end else begin
		if (wer2_is_error) begin
			wer2_wer_counter <= (wer2_wer_counter + 1'd1);
		end
	end
	if (wer2_i) begin
		wer2_toggle_i <= (~wer2_toggle_i);
	end
	decoding2_output_de <= 1'd1;
	if ((decoding2_input == 10'd852)) begin
		decoding2_output_de <= 1'd0;
		decoding2_output_c <= 1'd0;
	end
	if ((decoding2_input == 8'd171)) begin
		decoding2_output_de <= 1'd0;
		decoding2_output_c <= 1'd1;
	end
	if ((decoding2_input == 9'd340)) begin
		decoding2_output_de <= 1'd0;
		decoding2_output_c <= 2'd2;
	end
	if ((decoding2_input == 10'd683)) begin
		decoding2_output_de <= 1'd0;
		decoding2_output_c <= 2'd3;
	end
	decoding2_output_d[0] <= (decoding2_input[0] ^ decoding2_input[9]);
	decoding2_output_d[1] <= ((decoding2_input[1] ^ decoding2_input[0]) ^ (~decoding2_input[8]));
	decoding2_output_d[2] <= ((decoding2_input[2] ^ decoding2_input[1]) ^ (~decoding2_input[8]));
	decoding2_output_d[3] <= ((decoding2_input[3] ^ decoding2_input[2]) ^ (~decoding2_input[8]));
	decoding2_output_d[4] <= ((decoding2_input[4] ^ decoding2_input[3]) ^ (~decoding2_input[8]));
	decoding2_output_d[5] <= ((decoding2_input[5] ^ decoding2_input[4]) ^ (~decoding2_input[8]));
	decoding2_output_d[6] <= ((decoding2_input[6] ^ decoding2_input[5]) ^ (~decoding2_input[8]));
	decoding2_output_d[7] <= ((decoding2_input[7] ^ decoding2_input[6]) ^ (~decoding2_input[8]));
	decoding2_valid_o <= decoding2_valid_i;
	if ((~chansync_valid_i)) begin
		chansync_chan_synced <= 1'd0;
	end else begin
		if (chansync_some_control) begin
			if (chansync_all_control) begin
				chansync_chan_synced <= 1'd1;
			end else begin
				chansync_chan_synced <= 1'd0;
			end
		end
	end
	chansync_syncbuffer0_produce <= (chansync_syncbuffer0_produce + 1'd1);
	if (chansync_syncbuffer0_re) begin
		chansync_syncbuffer0_consume <= (chansync_syncbuffer0_consume + 1'd1);
	end
	chansync_syncbuffer1_produce <= (chansync_syncbuffer1_produce + 1'd1);
	if (chansync_syncbuffer1_re) begin
		chansync_syncbuffer1_consume <= (chansync_syncbuffer1_consume + 1'd1);
	end
	chansync_syncbuffer2_produce <= (chansync_syncbuffer2_produce + 1'd1);
	if (chansync_syncbuffer2_re) begin
		chansync_syncbuffer2_consume <= (chansync_syncbuffer2_consume + 1'd1);
	end
	syncpol_valid_o <= syncpol_valid_i;
	syncpol_r <= syncpol_data_in2_d;
	syncpol_g <= syncpol_data_in1_d;
	syncpol_b <= syncpol_data_in0_d;
	syncpol_de_r <= syncpol_data_in0_de;
	if ((syncpol_de_r & (~syncpol_data_in0_de))) begin
		syncpol_c_polarity <= syncpol_data_in0_c;
		syncpol_c_out <= 1'd0;
	end else begin
		syncpol_c_out <= (syncpol_data_in0_c ^ syncpol_c_polarity);
	end
	resdetection_de_r <= resdetection_de;
	if ((resdetection_valid_i & resdetection_de)) begin
		resdetection_hcounter <= (resdetection_hcounter + 1'd1);
	end else begin
		resdetection_hcounter <= 1'd0;
	end
	if (resdetection_valid_i) begin
		if (resdetection_pn_de) begin
			resdetection_hcounter_st <= resdetection_hcounter;
		end
	end else begin
		resdetection_hcounter_st <= 1'd0;
	end
	resdetection_vsync_r <= resdetection_vsync;
	if ((resdetection_valid_i & resdetection_p_vsync)) begin
		resdetection_vcounter <= 1'd0;
	end else begin
		if (resdetection_pn_de) begin
			resdetection_vcounter <= (resdetection_vcounter + 1'd1);
		end
	end
	if (resdetection_valid_i) begin
		if (resdetection_p_vsync) begin
			resdetection_vcounter_st <= resdetection_vcounter;
		end
	end else begin
		resdetection_vcounter_st <= 1'd0;
	end
	frame_de_r <= frame_de;
	frame_next_de0 <= frame_de;
	frame_next_vsync0 <= frame_vsync;
	frame_next_de1 <= frame_next_de0;
	frame_next_vsync1 <= frame_next_vsync0;
	frame_next_de2 <= frame_next_de1;
	frame_next_vsync2 <= frame_next_vsync1;
	frame_next_de3 <= frame_next_de2;
	frame_next_vsync3 <= frame_next_vsync2;
	frame_next_de4 <= frame_next_de3;
	frame_next_vsync4 <= frame_next_vsync3;
	frame_next_de5 <= frame_next_de4;
	frame_next_vsync5 <= frame_next_vsync4;
	frame_next_de6 <= frame_next_de5;
	frame_next_vsync6 <= frame_next_vsync5;
	frame_next_de7 <= frame_next_de6;
	frame_next_vsync7 <= frame_next_vsync6;
	frame_next_de8 <= frame_next_de7;
	frame_next_vsync8 <= frame_next_vsync7;
	frame_next_de9 <= frame_next_de8;
	frame_next_vsync9 <= frame_next_vsync8;
	frame_next_de10 <= frame_next_de9;
	frame_next_vsync10 <= frame_next_vsync9;
	frame_vsync_r <= frame_next_vsync10;
	frame_cur_word_valid <= 1'd0;
	if (frame_new_frame) begin
		frame_cur_word_valid <= (frame_pack_counter == 3'd7);
		frame_pack_counter <= 1'd0;
	end else begin
		if ((frame_chroma_downsampler_source_valid & frame_next_de10)) begin
			if ((frame_pack_counter == 3'd7)) begin
				frame_cur_word[15:0] <= frame_encoded_pixel;
			end
			if ((frame_pack_counter == 3'd6)) begin
				frame_cur_word[31:16] <= frame_encoded_pixel;
			end
			if ((frame_pack_counter == 3'd5)) begin
				frame_cur_word[47:32] <= frame_encoded_pixel;
			end
			if ((frame_pack_counter == 3'd4)) begin
				frame_cur_word[63:48] <= frame_encoded_pixel;
			end
			if ((frame_pack_counter == 2'd3)) begin
				frame_cur_word[79:64] <= frame_encoded_pixel;
			end
			if ((frame_pack_counter == 2'd2)) begin
				frame_cur_word[95:80] <= frame_encoded_pixel;
			end
			if ((frame_pack_counter == 1'd1)) begin
				frame_cur_word[111:96] <= frame_encoded_pixel;
			end
			if ((frame_pack_counter == 1'd0)) begin
				frame_cur_word[127:112] <= frame_encoded_pixel;
			end
			frame_cur_word_valid <= (frame_pack_counter == 3'd7);
			frame_pack_counter <= (frame_pack_counter + 1'd1);
		end
	end
	if (frame_new_frame) begin
		frame_fifo_sink_payload_sof <= 1'd1;
	end else begin
		if (frame_cur_word_valid) begin
			frame_fifo_sink_payload_sof <= 1'd0;
		end
	end
	if ((frame_fifo_sink_valid & (~frame_fifo_sink_ready))) begin
		frame_pix_overflow <= 1'd1;
	end else begin
		if (frame_pix_overflow_reset) begin
			frame_pix_overflow <= 1'd0;
		end
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n0 <= frame_rgb2ycbcr_sink_valid;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n1 <= frame_rgb2ycbcr_valid_n0;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n2 <= frame_rgb2ycbcr_valid_n1;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n3 <= frame_rgb2ycbcr_valid_n2;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n4 <= frame_rgb2ycbcr_valid_n3;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n5 <= frame_rgb2ycbcr_valid_n4;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n6 <= frame_rgb2ycbcr_valid_n5;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_valid_n7 <= frame_rgb2ycbcr_valid_n6;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n0 <= (frame_rgb2ycbcr_sink_valid & frame_rgb2ycbcr_sink_first);
		frame_rgb2ycbcr_last_n0 <= (frame_rgb2ycbcr_sink_valid & frame_rgb2ycbcr_sink_last);
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n1 <= frame_rgb2ycbcr_first_n0;
		frame_rgb2ycbcr_last_n1 <= frame_rgb2ycbcr_last_n0;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n2 <= frame_rgb2ycbcr_first_n1;
		frame_rgb2ycbcr_last_n2 <= frame_rgb2ycbcr_last_n1;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n3 <= frame_rgb2ycbcr_first_n2;
		frame_rgb2ycbcr_last_n3 <= frame_rgb2ycbcr_last_n2;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n4 <= frame_rgb2ycbcr_first_n3;
		frame_rgb2ycbcr_last_n4 <= frame_rgb2ycbcr_last_n3;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n5 <= frame_rgb2ycbcr_first_n4;
		frame_rgb2ycbcr_last_n5 <= frame_rgb2ycbcr_last_n4;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n6 <= frame_rgb2ycbcr_first_n5;
		frame_rgb2ycbcr_last_n6 <= frame_rgb2ycbcr_last_n5;
	end
	if (frame_rgb2ycbcr_pipe_ce) begin
		frame_rgb2ycbcr_first_n7 <= frame_rgb2ycbcr_first_n6;
		frame_rgb2ycbcr_last_n7 <= frame_rgb2ycbcr_last_n6;
	end
	if (frame_rgb2ycbcr_ce) begin
		frame_rgb2ycbcr_record0_rgb_n_r <= frame_rgb2ycbcr_sink_r;
		frame_rgb2ycbcr_record0_rgb_n_g <= frame_rgb2ycbcr_sink_g;
		frame_rgb2ycbcr_record0_rgb_n_b <= frame_rgb2ycbcr_sink_b;
		frame_rgb2ycbcr_record1_rgb_n_r <= frame_rgb2ycbcr_record0_rgb_n_r;
		frame_rgb2ycbcr_record1_rgb_n_g <= frame_rgb2ycbcr_record0_rgb_n_g;
		frame_rgb2ycbcr_record1_rgb_n_b <= frame_rgb2ycbcr_record0_rgb_n_b;
		frame_rgb2ycbcr_record2_rgb_n_r <= frame_rgb2ycbcr_record1_rgb_n_r;
		frame_rgb2ycbcr_record2_rgb_n_g <= frame_rgb2ycbcr_record1_rgb_n_g;
		frame_rgb2ycbcr_record2_rgb_n_b <= frame_rgb2ycbcr_record1_rgb_n_b;
		frame_rgb2ycbcr_record3_rgb_n_r <= frame_rgb2ycbcr_record2_rgb_n_r;
		frame_rgb2ycbcr_record3_rgb_n_g <= frame_rgb2ycbcr_record2_rgb_n_g;
		frame_rgb2ycbcr_record3_rgb_n_b <= frame_rgb2ycbcr_record2_rgb_n_b;
		frame_rgb2ycbcr_record4_rgb_n_r <= frame_rgb2ycbcr_record3_rgb_n_r;
		frame_rgb2ycbcr_record4_rgb_n_g <= frame_rgb2ycbcr_record3_rgb_n_g;
		frame_rgb2ycbcr_record4_rgb_n_b <= frame_rgb2ycbcr_record3_rgb_n_b;
		frame_rgb2ycbcr_record5_rgb_n_r <= frame_rgb2ycbcr_record4_rgb_n_r;
		frame_rgb2ycbcr_record5_rgb_n_g <= frame_rgb2ycbcr_record4_rgb_n_g;
		frame_rgb2ycbcr_record5_rgb_n_b <= frame_rgb2ycbcr_record4_rgb_n_b;
		frame_rgb2ycbcr_record6_rgb_n_r <= frame_rgb2ycbcr_record5_rgb_n_r;
		frame_rgb2ycbcr_record6_rgb_n_g <= frame_rgb2ycbcr_record5_rgb_n_g;
		frame_rgb2ycbcr_record6_rgb_n_b <= frame_rgb2ycbcr_record5_rgb_n_b;
		frame_rgb2ycbcr_record7_rgb_n_r <= frame_rgb2ycbcr_record6_rgb_n_r;
		frame_rgb2ycbcr_record7_rgb_n_g <= frame_rgb2ycbcr_record6_rgb_n_g;
		frame_rgb2ycbcr_record7_rgb_n_b <= frame_rgb2ycbcr_record6_rgb_n_b;
		frame_rgb2ycbcr_r_minus_g <= (frame_rgb2ycbcr_sink_r - frame_rgb2ycbcr_sink_g);
		frame_rgb2ycbcr_b_minus_g <= (frame_rgb2ycbcr_sink_b - frame_rgb2ycbcr_sink_g);
		frame_rgb2ycbcr_ca_mult_rg <= (frame_rgb2ycbcr_r_minus_g * $signed({1'd0, 6'd46}));
		frame_rgb2ycbcr_cb_mult_bg <= (frame_rgb2ycbcr_b_minus_g * $signed({1'd0, 4'd15}));
		frame_rgb2ycbcr_carg_plus_cbbg <= (frame_rgb2ycbcr_ca_mult_rg + frame_rgb2ycbcr_cb_mult_bg);
		frame_rgb2ycbcr_yraw <= (frame_rgb2ycbcr_carg_plus_cbbg[24:8] + $signed({1'd0, frame_rgb2ycbcr_record2_rgb_n_g}));
		frame_rgb2ycbcr_b_minus_yraw <= ($signed({1'd0, frame_rgb2ycbcr_record3_rgb_n_b}) - frame_rgb2ycbcr_yraw);
		frame_rgb2ycbcr_r_minus_yraw <= ($signed({1'd0, frame_rgb2ycbcr_record3_rgb_n_r}) - frame_rgb2ycbcr_yraw);
		frame_rgb2ycbcr_yraw_r0 <= frame_rgb2ycbcr_yraw;
		frame_rgb2ycbcr_cc_mult_ryraw <= (frame_rgb2ycbcr_b_minus_yraw * $signed({1'd0, 8'd141}));
		frame_rgb2ycbcr_cd_mult_byraw <= (frame_rgb2ycbcr_r_minus_yraw * $signed({1'd0, 8'd166}));
		frame_rgb2ycbcr_yraw_r1 <= frame_rgb2ycbcr_yraw_r0;
		frame_rgb2ycbcr_y <= (frame_rgb2ycbcr_yraw_r1 + $signed({1'd0, 5'd16}));
		frame_rgb2ycbcr_cb <= (frame_rgb2ycbcr_cc_mult_ryraw[19:8] + $signed({1'd0, 8'd128}));
		frame_rgb2ycbcr_cr <= (frame_rgb2ycbcr_cd_mult_byraw[19:8] + $signed({1'd0, 8'd128}));
		if ((frame_rgb2ycbcr_y > $signed({1'd0, 8'd255}))) begin
			frame_rgb2ycbcr_source_y <= 8'd255;
		end else begin
			if ((frame_rgb2ycbcr_y < $signed({1'd0, 1'd0}))) begin
				frame_rgb2ycbcr_source_y <= 1'd0;
			end else begin
				frame_rgb2ycbcr_source_y <= frame_rgb2ycbcr_y;
			end
		end
		if ((frame_rgb2ycbcr_cb > $signed({1'd0, 8'd255}))) begin
			frame_rgb2ycbcr_source_cb <= 8'd255;
		end else begin
			if ((frame_rgb2ycbcr_cb < $signed({1'd0, 1'd0}))) begin
				frame_rgb2ycbcr_source_cb <= 1'd0;
			end else begin
				frame_rgb2ycbcr_source_cb <= frame_rgb2ycbcr_cb;
			end
		end
		if ((frame_rgb2ycbcr_cr > $signed({1'd0, 8'd255}))) begin
			frame_rgb2ycbcr_source_cr <= 8'd255;
		end else begin
			if ((frame_rgb2ycbcr_cr < $signed({1'd0, 1'd0}))) begin
				frame_rgb2ycbcr_source_cr <= 1'd0;
			end else begin
				frame_rgb2ycbcr_source_cr <= frame_rgb2ycbcr_cr;
			end
		end
	end
	if (frame_chroma_downsampler_pipe_ce) begin
		frame_chroma_downsampler_valid_n0 <= frame_chroma_downsampler_sink_valid;
	end
	if (frame_chroma_downsampler_pipe_ce) begin
		frame_chroma_downsampler_valid_n1 <= frame_chroma_downsampler_valid_n0;
	end
	if (frame_chroma_downsampler_pipe_ce) begin
		frame_chroma_downsampler_valid_n2 <= frame_chroma_downsampler_valid_n1;
	end
	if (frame_chroma_downsampler_pipe_ce) begin
		frame_chroma_downsampler_first_n0 <= (frame_chroma_downsampler_sink_valid & frame_chroma_downsampler_sink_first);
		frame_chroma_downsampler_last_n0 <= (frame_chroma_downsampler_sink_valid & frame_chroma_downsampler_sink_last);
	end
	if (frame_chroma_downsampler_pipe_ce) begin
		frame_chroma_downsampler_first_n1 <= frame_chroma_downsampler_first_n0;
		frame_chroma_downsampler_last_n1 <= frame_chroma_downsampler_last_n0;
	end
	if (frame_chroma_downsampler_pipe_ce) begin
		frame_chroma_downsampler_first_n2 <= frame_chroma_downsampler_first_n1;
		frame_chroma_downsampler_last_n2 <= frame_chroma_downsampler_last_n1;
	end
	if (frame_chroma_downsampler_ce) begin
		frame_chroma_downsampler_record0_ycbcr_n_y <= frame_chroma_downsampler_sink_y;
		frame_chroma_downsampler_record0_ycbcr_n_cb <= frame_chroma_downsampler_sink_cb;
		frame_chroma_downsampler_record0_ycbcr_n_cr <= frame_chroma_downsampler_sink_cr;
		frame_chroma_downsampler_record1_ycbcr_n_y <= frame_chroma_downsampler_record0_ycbcr_n_y;
		frame_chroma_downsampler_record1_ycbcr_n_cb <= frame_chroma_downsampler_record0_ycbcr_n_cb;
		frame_chroma_downsampler_record1_ycbcr_n_cr <= frame_chroma_downsampler_record0_ycbcr_n_cr;
		frame_chroma_downsampler_record2_ycbcr_n_y <= frame_chroma_downsampler_record1_ycbcr_n_y;
		frame_chroma_downsampler_record2_ycbcr_n_cb <= frame_chroma_downsampler_record1_ycbcr_n_cb;
		frame_chroma_downsampler_record2_ycbcr_n_cr <= frame_chroma_downsampler_record1_ycbcr_n_cr;
		if ((frame_chroma_downsampler_first | (~frame_chroma_downsampler_parity))) begin
			frame_chroma_downsampler_parity <= 1'd1;
		end else begin
			frame_chroma_downsampler_parity <= 1'd0;
		end
		if (frame_chroma_downsampler_parity) begin
			frame_chroma_downsampler_cb_sum <= (frame_chroma_downsampler_sink_cb + frame_chroma_downsampler_record0_ycbcr_n_cb);
			frame_chroma_downsampler_cr_sum <= (frame_chroma_downsampler_sink_cr + frame_chroma_downsampler_record0_ycbcr_n_cr);
		end
		if (frame_chroma_downsampler_parity) begin
			frame_chroma_downsampler_source_y <= frame_chroma_downsampler_record1_ycbcr_n_y;
			frame_chroma_downsampler_source_cb_cr <= frame_chroma_downsampler_cr_mean;
		end else begin
			frame_chroma_downsampler_source_y <= frame_chroma_downsampler_record1_ycbcr_n_y;
			frame_chroma_downsampler_source_cb_cr <= frame_chroma_downsampler_cb_mean;
		end
	end
	frame_fifo_graycounter0_q_binary <= frame_fifo_graycounter0_q_next_binary;
	frame_fifo_graycounter0_q <= frame_fifo_graycounter0_q_next;
	frame_overflow_reset_toggle_o_r <= frame_overflow_reset_toggle_o;
	if (frame_overflow_reset_ack_i) begin
		frame_overflow_reset_ack_toggle_i <= (~frame_overflow_reset_ack_toggle_i);
	end
	if (hdmi_in0_pix_rst) begin
		charsync0_synced <= 1'd0;
		charsync0_data <= 10'd0;
		charsync0_raw_data1 <= 10'd0;
		charsync0_found_control <= 1'd0;
		charsync0_control_position <= 4'd0;
		charsync0_control_counter <= 3'd0;
		charsync0_previous_control_position <= 4'd0;
		charsync0_word_sel <= 4'd0;
		wer0_data_r <= 9'd0;
		wer0_transition_count <= 4'd0;
		wer0_is_control <= 1'd0;
		wer0_is_error <= 1'd0;
		wer0_period_counter <= 24'd0;
		wer0_period_done <= 1'd0;
		wer0_wer_counter <= 24'd0;
		wer0_wer_counter_r <= 24'd0;
		wer0_wer_counter_r_updated <= 1'd0;
		decoding0_valid_o <= 1'd0;
		decoding0_output_d <= 8'd0;
		decoding0_output_c <= 2'd0;
		decoding0_output_de <= 1'd0;
		charsync1_synced <= 1'd0;
		charsync1_data <= 10'd0;
		charsync1_raw_data1 <= 10'd0;
		charsync1_found_control <= 1'd0;
		charsync1_control_position <= 4'd0;
		charsync1_control_counter <= 3'd0;
		charsync1_previous_control_position <= 4'd0;
		charsync1_word_sel <= 4'd0;
		wer1_data_r <= 9'd0;
		wer1_transition_count <= 4'd0;
		wer1_is_control <= 1'd0;
		wer1_is_error <= 1'd0;
		wer1_period_counter <= 24'd0;
		wer1_period_done <= 1'd0;
		wer1_wer_counter <= 24'd0;
		wer1_wer_counter_r <= 24'd0;
		wer1_wer_counter_r_updated <= 1'd0;
		decoding1_valid_o <= 1'd0;
		decoding1_output_d <= 8'd0;
		decoding1_output_c <= 2'd0;
		decoding1_output_de <= 1'd0;
		charsync2_synced <= 1'd0;
		charsync2_data <= 10'd0;
		charsync2_raw_data1 <= 10'd0;
		charsync2_found_control <= 1'd0;
		charsync2_control_position <= 4'd0;
		charsync2_control_counter <= 3'd0;
		charsync2_previous_control_position <= 4'd0;
		charsync2_word_sel <= 4'd0;
		wer2_data_r <= 9'd0;
		wer2_transition_count <= 4'd0;
		wer2_is_control <= 1'd0;
		wer2_is_error <= 1'd0;
		wer2_period_counter <= 24'd0;
		wer2_period_done <= 1'd0;
		wer2_wer_counter <= 24'd0;
		wer2_wer_counter_r <= 24'd0;
		wer2_wer_counter_r_updated <= 1'd0;
		decoding2_valid_o <= 1'd0;
		decoding2_output_d <= 8'd0;
		decoding2_output_c <= 2'd0;
		decoding2_output_de <= 1'd0;
		chansync_chan_synced <= 1'd0;
		chansync_syncbuffer0_produce <= 3'd0;
		chansync_syncbuffer0_consume <= 3'd0;
		chansync_syncbuffer1_produce <= 3'd0;
		chansync_syncbuffer1_consume <= 3'd0;
		chansync_syncbuffer2_produce <= 3'd0;
		chansync_syncbuffer2_consume <= 3'd0;
		syncpol_valid_o <= 1'd0;
		syncpol_r <= 8'd0;
		syncpol_g <= 8'd0;
		syncpol_b <= 8'd0;
		syncpol_de_r <= 1'd0;
		syncpol_c_polarity <= 2'd0;
		syncpol_c_out <= 2'd0;
		resdetection_de_r <= 1'd0;
		resdetection_hcounter <= 11'd0;
		resdetection_hcounter_st <= 11'd0;
		resdetection_vsync_r <= 1'd0;
		resdetection_vcounter <= 11'd0;
		resdetection_vcounter_st <= 11'd0;
		frame_de_r <= 1'd0;
		frame_rgb2ycbcr_source_y <= 8'd0;
		frame_rgb2ycbcr_source_cb <= 8'd0;
		frame_rgb2ycbcr_source_cr <= 8'd0;
		frame_rgb2ycbcr_record0_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record0_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record0_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_record1_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record1_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record1_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_record2_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record2_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record2_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_record3_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record3_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record3_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_record4_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record4_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record4_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_record5_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record5_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record5_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_record6_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record6_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record6_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_record7_rgb_n_r <= 8'd0;
		frame_rgb2ycbcr_record7_rgb_n_g <= 8'd0;
		frame_rgb2ycbcr_record7_rgb_n_b <= 8'd0;
		frame_rgb2ycbcr_r_minus_g <= 9'sd512;
		frame_rgb2ycbcr_b_minus_g <= 9'sd512;
		frame_rgb2ycbcr_ca_mult_rg <= 17'sd131072;
		frame_rgb2ycbcr_cb_mult_bg <= 17'sd131072;
		frame_rgb2ycbcr_carg_plus_cbbg <= 25'sd33554432;
		frame_rgb2ycbcr_yraw <= 11'sd2048;
		frame_rgb2ycbcr_b_minus_yraw <= 12'sd4096;
		frame_rgb2ycbcr_r_minus_yraw <= 12'sd4096;
		frame_rgb2ycbcr_yraw_r0 <= 11'sd2048;
		frame_rgb2ycbcr_cc_mult_ryraw <= 20'sd1048576;
		frame_rgb2ycbcr_cd_mult_byraw <= 20'sd1048576;
		frame_rgb2ycbcr_yraw_r1 <= 11'sd2048;
		frame_rgb2ycbcr_y <= 11'sd2048;
		frame_rgb2ycbcr_cb <= 12'sd4096;
		frame_rgb2ycbcr_cr <= 12'sd4096;
		frame_rgb2ycbcr_valid_n0 <= 1'd0;
		frame_rgb2ycbcr_valid_n1 <= 1'd0;
		frame_rgb2ycbcr_valid_n2 <= 1'd0;
		frame_rgb2ycbcr_valid_n3 <= 1'd0;
		frame_rgb2ycbcr_valid_n4 <= 1'd0;
		frame_rgb2ycbcr_valid_n5 <= 1'd0;
		frame_rgb2ycbcr_valid_n6 <= 1'd0;
		frame_rgb2ycbcr_valid_n7 <= 1'd0;
		frame_rgb2ycbcr_first_n0 <= 1'd0;
		frame_rgb2ycbcr_last_n0 <= 1'd0;
		frame_rgb2ycbcr_first_n1 <= 1'd0;
		frame_rgb2ycbcr_last_n1 <= 1'd0;
		frame_rgb2ycbcr_first_n2 <= 1'd0;
		frame_rgb2ycbcr_last_n2 <= 1'd0;
		frame_rgb2ycbcr_first_n3 <= 1'd0;
		frame_rgb2ycbcr_last_n3 <= 1'd0;
		frame_rgb2ycbcr_first_n4 <= 1'd0;
		frame_rgb2ycbcr_last_n4 <= 1'd0;
		frame_rgb2ycbcr_first_n5 <= 1'd0;
		frame_rgb2ycbcr_last_n5 <= 1'd0;
		frame_rgb2ycbcr_first_n6 <= 1'd0;
		frame_rgb2ycbcr_last_n6 <= 1'd0;
		frame_rgb2ycbcr_first_n7 <= 1'd0;
		frame_rgb2ycbcr_last_n7 <= 1'd0;
		frame_chroma_downsampler_source_y <= 8'd0;
		frame_chroma_downsampler_source_cb_cr <= 8'd0;
		frame_chroma_downsampler_record0_ycbcr_n_y <= 8'd0;
		frame_chroma_downsampler_record0_ycbcr_n_cb <= 8'd0;
		frame_chroma_downsampler_record0_ycbcr_n_cr <= 8'd0;
		frame_chroma_downsampler_record1_ycbcr_n_y <= 8'd0;
		frame_chroma_downsampler_record1_ycbcr_n_cb <= 8'd0;
		frame_chroma_downsampler_record1_ycbcr_n_cr <= 8'd0;
		frame_chroma_downsampler_record2_ycbcr_n_y <= 8'd0;
		frame_chroma_downsampler_record2_ycbcr_n_cb <= 8'd0;
		frame_chroma_downsampler_record2_ycbcr_n_cr <= 8'd0;
		frame_chroma_downsampler_parity <= 1'd0;
		frame_chroma_downsampler_cb_sum <= 9'd0;
		frame_chroma_downsampler_cr_sum <= 9'd0;
		frame_chroma_downsampler_valid_n0 <= 1'd0;
		frame_chroma_downsampler_valid_n1 <= 1'd0;
		frame_chroma_downsampler_valid_n2 <= 1'd0;
		frame_chroma_downsampler_first_n0 <= 1'd0;
		frame_chroma_downsampler_last_n0 <= 1'd0;
		frame_chroma_downsampler_first_n1 <= 1'd0;
		frame_chroma_downsampler_last_n1 <= 1'd0;
		frame_chroma_downsampler_first_n2 <= 1'd0;
		frame_chroma_downsampler_last_n2 <= 1'd0;
		frame_next_de0 <= 1'd0;
		frame_next_vsync0 <= 1'd0;
		frame_next_de1 <= 1'd0;
		frame_next_vsync1 <= 1'd0;
		frame_next_de2 <= 1'd0;
		frame_next_vsync2 <= 1'd0;
		frame_next_de3 <= 1'd0;
		frame_next_vsync3 <= 1'd0;
		frame_next_de4 <= 1'd0;
		frame_next_vsync4 <= 1'd0;
		frame_next_de5 <= 1'd0;
		frame_next_vsync5 <= 1'd0;
		frame_next_de6 <= 1'd0;
		frame_next_vsync6 <= 1'd0;
		frame_next_de7 <= 1'd0;
		frame_next_vsync7 <= 1'd0;
		frame_next_de8 <= 1'd0;
		frame_next_vsync8 <= 1'd0;
		frame_next_de9 <= 1'd0;
		frame_next_vsync9 <= 1'd0;
		frame_next_de10 <= 1'd0;
		frame_next_vsync10 <= 1'd0;
		frame_vsync_r <= 1'd0;
		frame_cur_word <= 128'd0;
		frame_cur_word_valid <= 1'd0;
		frame_pack_counter <= 3'd0;
		frame_fifo_graycounter0_q <= 10'd0;
		frame_fifo_graycounter0_q_binary <= 10'd0;
		frame_pix_overflow <= 1'd0;
	end
	xilinxmultiregimpl45_regs0 <= frame_fifo_graycounter1_q;
	xilinxmultiregimpl45_regs1 <= xilinxmultiregimpl45_regs0;
	xilinxmultiregimpl47_regs0 <= frame_overflow_reset_toggle_i;
	xilinxmultiregimpl47_regs1 <= xilinxmultiregimpl47_regs0;
end

always @(posedge hdmi_out0_pix_clk) begin
	hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary <= hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary;
	hdmi_out0_dram_port_cmd_fifo_graycounter0_q <= hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next;
	hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary <= hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary;
	hdmi_out0_dram_port_rdata_fifo_graycounter1_q <= hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next;
	if (hdmi_out0_dram_port_counter_ce) begin
		hdmi_out0_dram_port_counter <= (hdmi_out0_dram_port_counter + 1'd1);
	end
	if ((hdmi_out0_dram_port_rdata_converter_source_valid & hdmi_out0_dram_port_rdata_converter_source_ready)) begin
		hdmi_out0_dram_port_rdata_chunk <= {hdmi_out0_dram_port_rdata_chunk[6:0], hdmi_out0_dram_port_rdata_chunk[7]};
	end
	if (((hdmi_out0_dram_port_cmd_buffer_syncfifo_we & hdmi_out0_dram_port_cmd_buffer_syncfifo_writable) & (~hdmi_out0_dram_port_cmd_buffer_replace))) begin
		hdmi_out0_dram_port_cmd_buffer_produce <= (hdmi_out0_dram_port_cmd_buffer_produce + 1'd1);
	end
	if (hdmi_out0_dram_port_cmd_buffer_do_read) begin
		hdmi_out0_dram_port_cmd_buffer_consume <= (hdmi_out0_dram_port_cmd_buffer_consume + 1'd1);
	end
	if (((hdmi_out0_dram_port_cmd_buffer_syncfifo_we & hdmi_out0_dram_port_cmd_buffer_syncfifo_writable) & (~hdmi_out0_dram_port_cmd_buffer_replace))) begin
		if ((~hdmi_out0_dram_port_cmd_buffer_do_read)) begin
			hdmi_out0_dram_port_cmd_buffer_level <= (hdmi_out0_dram_port_cmd_buffer_level + 1'd1);
		end
	end else begin
		if (hdmi_out0_dram_port_cmd_buffer_do_read) begin
			hdmi_out0_dram_port_cmd_buffer_level <= (hdmi_out0_dram_port_cmd_buffer_level - 1'd1);
		end
	end
	if (hdmi_out0_dram_port_rdata_buffer_pipe_ce) begin
		hdmi_out0_dram_port_rdata_buffer_valid_n <= hdmi_out0_dram_port_rdata_buffer_sink_valid;
	end
	if (hdmi_out0_dram_port_rdata_buffer_pipe_ce) begin
		hdmi_out0_dram_port_rdata_buffer_first_n <= (hdmi_out0_dram_port_rdata_buffer_sink_valid & hdmi_out0_dram_port_rdata_buffer_sink_first);
		hdmi_out0_dram_port_rdata_buffer_last_n <= (hdmi_out0_dram_port_rdata_buffer_sink_valid & hdmi_out0_dram_port_rdata_buffer_sink_last);
	end
	if (hdmi_out0_dram_port_rdata_buffer_pipe_ce) begin
		hdmi_out0_dram_port_rdata_buffer_source_payload_data <= hdmi_out0_dram_port_rdata_buffer_sink_payload_data;
	end
	if ((hdmi_out0_dram_port_rdata_converter_converter_source_valid & hdmi_out0_dram_port_rdata_converter_converter_source_ready)) begin
		if (hdmi_out0_dram_port_rdata_converter_converter_last) begin
			hdmi_out0_dram_port_rdata_converter_converter_mux <= 1'd0;
		end else begin
			hdmi_out0_dram_port_rdata_converter_converter_mux <= (hdmi_out0_dram_port_rdata_converter_converter_mux + 1'd1);
		end
	end
	hdmi_out0_de_r <= hdmi_out0_core_source_source_param_de;
	hdmi_out0_core_source_valid_d <= hdmi_out0_core_source_source_valid;
	hdmi_out0_core_source_data_d <= hdmi_out0_core_source_source_payload_data;
	if (hdmi_out0_core_underflow_enable) begin
		if ((~hdmi_out0_core_source_source_valid)) begin
			hdmi_out0_core_underflow_counter <= (hdmi_out0_core_underflow_counter + 1'd1);
		end
	end else begin
		hdmi_out0_core_underflow_counter <= 1'd0;
	end
	if (hdmi_out0_core_underflow_update) begin
		hdmi_out0_core_underflow_counter_status <= hdmi_out0_core_underflow_counter;
	end
	hdmi_out0_core_initiator_cdc_graycounter1_q_binary <= hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary;
	hdmi_out0_core_initiator_cdc_graycounter1_q <= hdmi_out0_core_initiator_cdc_graycounter1_q_next;
	if ((~hdmi_out0_core_timinggenerator_sink_valid)) begin
		hdmi_out0_core_timinggenerator_hactive <= 1'd0;
		hdmi_out0_core_timinggenerator_vactive <= 1'd0;
		hdmi_out0_core_timinggenerator_hcounter <= 1'd0;
		hdmi_out0_core_timinggenerator_vcounter <= 1'd0;
	end else begin
		if (hdmi_out0_core_timinggenerator_source_ready) begin
			hdmi_out0_core_timinggenerator_source_last <= 1'd0;
			hdmi_out0_core_timinggenerator_hcounter <= (hdmi_out0_core_timinggenerator_hcounter + 1'd1);
			if ((hdmi_out0_core_timinggenerator_hcounter == 1'd0)) begin
				hdmi_out0_core_timinggenerator_hactive <= 1'd1;
			end
			if ((hdmi_out0_core_timinggenerator_hcounter == hdmi_out0_core_timinggenerator_sink_payload_hres)) begin
				hdmi_out0_core_timinggenerator_hactive <= 1'd0;
			end
			if ((hdmi_out0_core_timinggenerator_hcounter == hdmi_out0_core_timinggenerator_sink_payload_hsync_start)) begin
				hdmi_out0_core_timinggenerator_source_payload_hsync <= 1'd1;
			end
			if ((hdmi_out0_core_timinggenerator_hcounter == hdmi_out0_core_timinggenerator_sink_payload_hsync_end)) begin
				hdmi_out0_core_timinggenerator_source_payload_hsync <= 1'd0;
			end
			if ((hdmi_out0_core_timinggenerator_hcounter == hdmi_out0_core_timinggenerator_sink_payload_hscan)) begin
				hdmi_out0_core_timinggenerator_hcounter <= 1'd0;
				if ((hdmi_out0_core_timinggenerator_vcounter == hdmi_out0_core_timinggenerator_sink_payload_vscan)) begin
					hdmi_out0_core_timinggenerator_vcounter <= 1'd0;
					hdmi_out0_core_timinggenerator_source_last <= 1'd1;
				end else begin
					hdmi_out0_core_timinggenerator_vcounter <= (hdmi_out0_core_timinggenerator_vcounter + 1'd1);
				end
			end
			if ((hdmi_out0_core_timinggenerator_vcounter == 1'd0)) begin
				hdmi_out0_core_timinggenerator_vactive <= 1'd1;
			end
			if ((hdmi_out0_core_timinggenerator_vcounter == hdmi_out0_core_timinggenerator_sink_payload_vres)) begin
				hdmi_out0_core_timinggenerator_vactive <= 1'd0;
			end
			if ((hdmi_out0_core_timinggenerator_vcounter == hdmi_out0_core_timinggenerator_sink_payload_vsync_start)) begin
				hdmi_out0_core_timinggenerator_source_payload_vsync <= 1'd1;
			end
			if ((hdmi_out0_core_timinggenerator_vcounter == hdmi_out0_core_timinggenerator_sink_payload_vsync_end)) begin
				hdmi_out0_core_timinggenerator_source_payload_vsync <= 1'd0;
			end
		end
	end
	if (hdmi_out0_core_dmareader_request_issued) begin
		if ((~hdmi_out0_core_dmareader_data_dequeued)) begin
			hdmi_out0_core_dmareader_rsv_level <= (hdmi_out0_core_dmareader_rsv_level + 1'd1);
		end
	end else begin
		if (hdmi_out0_core_dmareader_data_dequeued) begin
			hdmi_out0_core_dmareader_rsv_level <= (hdmi_out0_core_dmareader_rsv_level - 1'd1);
		end
	end
	if (hdmi_out0_core_dmareader_fifo_syncfifo_re) begin
		hdmi_out0_core_dmareader_fifo_readable <= 1'd1;
	end else begin
		if (hdmi_out0_core_dmareader_fifo_re) begin
			hdmi_out0_core_dmareader_fifo_readable <= 1'd0;
		end
	end
	if (((hdmi_out0_core_dmareader_fifo_syncfifo_we & hdmi_out0_core_dmareader_fifo_syncfifo_writable) & (~hdmi_out0_core_dmareader_fifo_replace))) begin
		hdmi_out0_core_dmareader_fifo_produce <= (hdmi_out0_core_dmareader_fifo_produce + 1'd1);
	end
	if (hdmi_out0_core_dmareader_fifo_do_read) begin
		hdmi_out0_core_dmareader_fifo_consume <= (hdmi_out0_core_dmareader_fifo_consume + 1'd1);
	end
	if (((hdmi_out0_core_dmareader_fifo_syncfifo_we & hdmi_out0_core_dmareader_fifo_syncfifo_writable) & (~hdmi_out0_core_dmareader_fifo_replace))) begin
		if ((~hdmi_out0_core_dmareader_fifo_do_read)) begin
			hdmi_out0_core_dmareader_fifo_level0 <= (hdmi_out0_core_dmareader_fifo_level0 + 1'd1);
		end
	end else begin
		if (hdmi_out0_core_dmareader_fifo_do_read) begin
			hdmi_out0_core_dmareader_fifo_level0 <= (hdmi_out0_core_dmareader_fifo_level0 - 1'd1);
		end
	end
	videoout_state <= videoout_next_state;
	if (hdmi_out0_core_dmareader_offset_videoout_next_value_ce) begin
		hdmi_out0_core_dmareader_offset <= hdmi_out0_core_dmareader_offset_videoout_next_value;
	end
	hdmi_out0_core_toggle_o_r <= hdmi_out0_core_toggle_o;
	if ((hdmi_out0_resetinserter_sink_sink_valid & hdmi_out0_resetinserter_sink_sink_ready)) begin
		hdmi_out0_resetinserter_parity_in <= (~hdmi_out0_resetinserter_parity_in);
	end
	if ((hdmi_out0_resetinserter_source_source_valid & hdmi_out0_resetinserter_source_source_ready)) begin
		hdmi_out0_resetinserter_parity_out <= (~hdmi_out0_resetinserter_parity_out);
	end
	if (((hdmi_out0_resetinserter_y_fifo_syncfifo_we & hdmi_out0_resetinserter_y_fifo_syncfifo_writable) & (~hdmi_out0_resetinserter_y_fifo_replace))) begin
		hdmi_out0_resetinserter_y_fifo_produce <= (hdmi_out0_resetinserter_y_fifo_produce + 1'd1);
	end
	if (hdmi_out0_resetinserter_y_fifo_do_read) begin
		hdmi_out0_resetinserter_y_fifo_consume <= (hdmi_out0_resetinserter_y_fifo_consume + 1'd1);
	end
	if (((hdmi_out0_resetinserter_y_fifo_syncfifo_we & hdmi_out0_resetinserter_y_fifo_syncfifo_writable) & (~hdmi_out0_resetinserter_y_fifo_replace))) begin
		if ((~hdmi_out0_resetinserter_y_fifo_do_read)) begin
			hdmi_out0_resetinserter_y_fifo_level <= (hdmi_out0_resetinserter_y_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi_out0_resetinserter_y_fifo_do_read) begin
			hdmi_out0_resetinserter_y_fifo_level <= (hdmi_out0_resetinserter_y_fifo_level - 1'd1);
		end
	end
	if (((hdmi_out0_resetinserter_cb_fifo_syncfifo_we & hdmi_out0_resetinserter_cb_fifo_syncfifo_writable) & (~hdmi_out0_resetinserter_cb_fifo_replace))) begin
		hdmi_out0_resetinserter_cb_fifo_produce <= (hdmi_out0_resetinserter_cb_fifo_produce + 1'd1);
	end
	if (hdmi_out0_resetinserter_cb_fifo_do_read) begin
		hdmi_out0_resetinserter_cb_fifo_consume <= (hdmi_out0_resetinserter_cb_fifo_consume + 1'd1);
	end
	if (((hdmi_out0_resetinserter_cb_fifo_syncfifo_we & hdmi_out0_resetinserter_cb_fifo_syncfifo_writable) & (~hdmi_out0_resetinserter_cb_fifo_replace))) begin
		if ((~hdmi_out0_resetinserter_cb_fifo_do_read)) begin
			hdmi_out0_resetinserter_cb_fifo_level <= (hdmi_out0_resetinserter_cb_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi_out0_resetinserter_cb_fifo_do_read) begin
			hdmi_out0_resetinserter_cb_fifo_level <= (hdmi_out0_resetinserter_cb_fifo_level - 1'd1);
		end
	end
	if (((hdmi_out0_resetinserter_cr_fifo_syncfifo_we & hdmi_out0_resetinserter_cr_fifo_syncfifo_writable) & (~hdmi_out0_resetinserter_cr_fifo_replace))) begin
		hdmi_out0_resetinserter_cr_fifo_produce <= (hdmi_out0_resetinserter_cr_fifo_produce + 1'd1);
	end
	if (hdmi_out0_resetinserter_cr_fifo_do_read) begin
		hdmi_out0_resetinserter_cr_fifo_consume <= (hdmi_out0_resetinserter_cr_fifo_consume + 1'd1);
	end
	if (((hdmi_out0_resetinserter_cr_fifo_syncfifo_we & hdmi_out0_resetinserter_cr_fifo_syncfifo_writable) & (~hdmi_out0_resetinserter_cr_fifo_replace))) begin
		if ((~hdmi_out0_resetinserter_cr_fifo_do_read)) begin
			hdmi_out0_resetinserter_cr_fifo_level <= (hdmi_out0_resetinserter_cr_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi_out0_resetinserter_cr_fifo_do_read) begin
			hdmi_out0_resetinserter_cr_fifo_level <= (hdmi_out0_resetinserter_cr_fifo_level - 1'd1);
		end
	end
	if (hdmi_out0_resetinserter_reset) begin
		hdmi_out0_resetinserter_y_fifo_level <= 3'd0;
		hdmi_out0_resetinserter_y_fifo_produce <= 2'd0;
		hdmi_out0_resetinserter_y_fifo_consume <= 2'd0;
		hdmi_out0_resetinserter_cb_fifo_level <= 3'd0;
		hdmi_out0_resetinserter_cb_fifo_produce <= 2'd0;
		hdmi_out0_resetinserter_cb_fifo_consume <= 2'd0;
		hdmi_out0_resetinserter_cr_fifo_level <= 3'd0;
		hdmi_out0_resetinserter_cr_fifo_produce <= 2'd0;
		hdmi_out0_resetinserter_cr_fifo_consume <= 2'd0;
		hdmi_out0_resetinserter_parity_in <= 1'd0;
		hdmi_out0_resetinserter_parity_out <= 1'd0;
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_valid_n0 <= hdmi_out0_sink_valid;
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_valid_n1 <= hdmi_out0_valid_n0;
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_valid_n2 <= hdmi_out0_valid_n1;
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_valid_n3 <= hdmi_out0_valid_n2;
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_first_n0 <= (hdmi_out0_sink_valid & hdmi_out0_sink_first);
		hdmi_out0_last_n0 <= (hdmi_out0_sink_valid & hdmi_out0_sink_last);
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_first_n1 <= hdmi_out0_first_n0;
		hdmi_out0_last_n1 <= hdmi_out0_last_n0;
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_first_n2 <= hdmi_out0_first_n1;
		hdmi_out0_last_n2 <= hdmi_out0_last_n1;
	end
	if (hdmi_out0_pipe_ce) begin
		hdmi_out0_first_n3 <= hdmi_out0_first_n2;
		hdmi_out0_last_n3 <= hdmi_out0_last_n2;
	end
	if (hdmi_out0_ce) begin
		hdmi_out0_record0_ycbcr_n_y <= hdmi_out0_sink_y;
		hdmi_out0_record0_ycbcr_n_cb <= hdmi_out0_sink_cb;
		hdmi_out0_record0_ycbcr_n_cr <= hdmi_out0_sink_cr;
		hdmi_out0_record1_ycbcr_n_y <= hdmi_out0_record0_ycbcr_n_y;
		hdmi_out0_record1_ycbcr_n_cb <= hdmi_out0_record0_ycbcr_n_cb;
		hdmi_out0_record1_ycbcr_n_cr <= hdmi_out0_record0_ycbcr_n_cr;
		hdmi_out0_record2_ycbcr_n_y <= hdmi_out0_record1_ycbcr_n_y;
		hdmi_out0_record2_ycbcr_n_cb <= hdmi_out0_record1_ycbcr_n_cb;
		hdmi_out0_record2_ycbcr_n_cr <= hdmi_out0_record1_ycbcr_n_cr;
		hdmi_out0_record3_ycbcr_n_y <= hdmi_out0_record2_ycbcr_n_y;
		hdmi_out0_record3_ycbcr_n_cb <= hdmi_out0_record2_ycbcr_n_cb;
		hdmi_out0_record3_ycbcr_n_cr <= hdmi_out0_record2_ycbcr_n_cr;
		hdmi_out0_cb_minus_coffset <= (hdmi_out0_sink_cb - 8'd128);
		hdmi_out0_cr_minus_coffset <= (hdmi_out0_sink_cr - 8'd128);
		hdmi_out0_y_minus_yoffset <= (hdmi_out0_record0_ycbcr_n_y - 5'd16);
		hdmi_out0_cr_minus_coffset_mult_acoef <= (hdmi_out0_cr_minus_coffset * $signed({1'd0, 7'd98}));
		hdmi_out0_cb_minus_coffset_mult_bcoef <= (hdmi_out0_cb_minus_coffset * 5'sd23);
		hdmi_out0_cr_minus_coffset_mult_ccoef <= (hdmi_out0_cr_minus_coffset * 6'sd41);
		hdmi_out0_cb_minus_coffset_mult_dcoef <= (hdmi_out0_cb_minus_coffset * $signed({1'd0, 7'd116}));
		hdmi_out0_r <= (hdmi_out0_y_minus_yoffset + hdmi_out0_cr_minus_coffset_mult_acoef[19:6]);
		hdmi_out0_g <= ((hdmi_out0_y_minus_yoffset + hdmi_out0_cb_minus_coffset_mult_bcoef[19:6]) + hdmi_out0_cr_minus_coffset_mult_ccoef[19:6]);
		hdmi_out0_b <= (hdmi_out0_y_minus_yoffset + hdmi_out0_cb_minus_coffset_mult_dcoef[19:6]);
		if ((hdmi_out0_r > $signed({1'd0, 8'd255}))) begin
			hdmi_out0_source_r <= 8'd255;
		end else begin
			if ((hdmi_out0_r < $signed({1'd0, 1'd0}))) begin
				hdmi_out0_source_r <= 1'd0;
			end else begin
				hdmi_out0_source_r <= hdmi_out0_r;
			end
		end
		if ((hdmi_out0_g > $signed({1'd0, 8'd255}))) begin
			hdmi_out0_source_g <= 8'd255;
		end else begin
			if ((hdmi_out0_g < $signed({1'd0, 1'd0}))) begin
				hdmi_out0_source_g <= 1'd0;
			end else begin
				hdmi_out0_source_g <= hdmi_out0_g;
			end
		end
		if ((hdmi_out0_b > $signed({1'd0, 8'd255}))) begin
			hdmi_out0_source_b <= 8'd255;
		end else begin
			if ((hdmi_out0_b < $signed({1'd0, 1'd0}))) begin
				hdmi_out0_source_b <= 1'd0;
			end else begin
				hdmi_out0_source_b <= hdmi_out0_b;
			end
		end
	end
	hdmi_out0_next_s0 <= hdmi_out0_sink_payload_hsync;
	hdmi_out0_next_s1 <= hdmi_out0_next_s0;
	hdmi_out0_next_s2 <= hdmi_out0_next_s1;
	hdmi_out0_next_s3 <= hdmi_out0_next_s2;
	hdmi_out0_next_s4 <= hdmi_out0_next_s3;
	hdmi_out0_next_s5 <= hdmi_out0_next_s4;
	hdmi_out0_next_s6 <= hdmi_out0_sink_payload_vsync;
	hdmi_out0_next_s7 <= hdmi_out0_next_s6;
	hdmi_out0_next_s8 <= hdmi_out0_next_s7;
	hdmi_out0_next_s9 <= hdmi_out0_next_s8;
	hdmi_out0_next_s10 <= hdmi_out0_next_s9;
	hdmi_out0_next_s11 <= hdmi_out0_next_s10;
	hdmi_out0_next_s12 <= hdmi_out0_sink_payload_de;
	hdmi_out0_next_s13 <= hdmi_out0_next_s12;
	hdmi_out0_next_s14 <= hdmi_out0_next_s13;
	hdmi_out0_next_s15 <= hdmi_out0_next_s14;
	hdmi_out0_next_s16 <= hdmi_out0_next_s15;
	hdmi_out0_next_s17 <= hdmi_out0_next_s16;
	hdmi_out0_driver_s7hdmioutclocking_ce <= (~hdmi_out0_pix_rst);
	hdmi_out0_driver_hdmi_phy_es0_ce <= (~hdmi_out0_pix_rst);
	hdmi_out0_driver_hdmi_phy_es0_n1d <= (((((((hdmi_out0_driver_hdmi_phy_es0_d0[0] + hdmi_out0_driver_hdmi_phy_es0_d0[1]) + hdmi_out0_driver_hdmi_phy_es0_d0[2]) + hdmi_out0_driver_hdmi_phy_es0_d0[3]) + hdmi_out0_driver_hdmi_phy_es0_d0[4]) + hdmi_out0_driver_hdmi_phy_es0_d0[5]) + hdmi_out0_driver_hdmi_phy_es0_d0[6]) + hdmi_out0_driver_hdmi_phy_es0_d0[7]);
	hdmi_out0_driver_hdmi_phy_es0_d1 <= hdmi_out0_driver_hdmi_phy_es0_d0;
	hdmi_out0_driver_hdmi_phy_es0_q_m[0] <= hdmi_out0_driver_hdmi_phy_es0_d1[0];
	hdmi_out0_driver_hdmi_phy_es0_q_m[1] <= ((hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_q_m[2] <= ((((hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_q_m[3] <= ((((((hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_q_m[4] <= ((((((((hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_q_m[5] <= ((((((((((hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_q_m[6] <= ((((((((((((hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[6]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_q_m[7] <= ((((((((((((((hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[6]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es0_d1[7]) ^ hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_q_m[8] <= (~hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es0_n0q_m <= ((((((((~hdmi_out0_driver_hdmi_phy_es0_q_m[0]) + (~hdmi_out0_driver_hdmi_phy_es0_q_m[1])) + (~hdmi_out0_driver_hdmi_phy_es0_q_m[2])) + (~hdmi_out0_driver_hdmi_phy_es0_q_m[3])) + (~hdmi_out0_driver_hdmi_phy_es0_q_m[4])) + (~hdmi_out0_driver_hdmi_phy_es0_q_m[5])) + (~hdmi_out0_driver_hdmi_phy_es0_q_m[6])) + (~hdmi_out0_driver_hdmi_phy_es0_q_m[7]));
	hdmi_out0_driver_hdmi_phy_es0_n1q_m <= (((((((hdmi_out0_driver_hdmi_phy_es0_q_m[0] + hdmi_out0_driver_hdmi_phy_es0_q_m[1]) + hdmi_out0_driver_hdmi_phy_es0_q_m[2]) + hdmi_out0_driver_hdmi_phy_es0_q_m[3]) + hdmi_out0_driver_hdmi_phy_es0_q_m[4]) + hdmi_out0_driver_hdmi_phy_es0_q_m[5]) + hdmi_out0_driver_hdmi_phy_es0_q_m[6]) + hdmi_out0_driver_hdmi_phy_es0_q_m[7]);
	hdmi_out0_driver_hdmi_phy_es0_q_m_r <= hdmi_out0_driver_hdmi_phy_es0_q_m;
	hdmi_out0_driver_hdmi_phy_es0_new_c0 <= hdmi_out0_driver_hdmi_phy_es0_c;
	hdmi_out0_driver_hdmi_phy_es0_new_de0 <= hdmi_out0_driver_hdmi_phy_es0_de;
	hdmi_out0_driver_hdmi_phy_es0_new_c1 <= hdmi_out0_driver_hdmi_phy_es0_new_c0;
	hdmi_out0_driver_hdmi_phy_es0_new_de1 <= hdmi_out0_driver_hdmi_phy_es0_new_de0;
	hdmi_out0_driver_hdmi_phy_es0_new_c2 <= hdmi_out0_driver_hdmi_phy_es0_new_c1;
	hdmi_out0_driver_hdmi_phy_es0_new_de2 <= hdmi_out0_driver_hdmi_phy_es0_new_de1;
	if (hdmi_out0_driver_hdmi_phy_es0_new_de2) begin
		if (((hdmi_out0_driver_hdmi_phy_es0_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es0_n1q_m == hdmi_out0_driver_hdmi_phy_es0_n0q_m)}))) begin
			hdmi_out0_driver_hdmi_phy_es0_out[9] <= (~hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]);
			hdmi_out0_driver_hdmi_phy_es0_out[8] <= hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
			if (hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]) begin
				hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0];
				hdmi_out0_driver_hdmi_phy_es0_cnt <= ((hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n0q_m}));
			end else begin
				hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= (~hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0]);
				hdmi_out0_driver_hdmi_phy_es0_cnt <= ((hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n1q_m}));
			end
		end else begin
			if ((((~hdmi_out0_driver_hdmi_phy_es0_cnt[5]) & $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es0_n1q_m > hdmi_out0_driver_hdmi_phy_es0_n0q_m)})) | (hdmi_out0_driver_hdmi_phy_es0_cnt[5] & $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es0_n0q_m > hdmi_out0_driver_hdmi_phy_es0_n1q_m)})))) begin
				hdmi_out0_driver_hdmi_phy_es0_out[9] <= 1'd1;
				hdmi_out0_driver_hdmi_phy_es0_out[8] <= hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
				hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= (~hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0]);
				hdmi_out0_driver_hdmi_phy_es0_cnt <= (((hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, {hdmi_out0_driver_hdmi_phy_es0_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n1q_m}));
			end else begin
				hdmi_out0_driver_hdmi_phy_es0_out[9] <= 1'd0;
				hdmi_out0_driver_hdmi_phy_es0_out[8] <= hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
				hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0];
				hdmi_out0_driver_hdmi_phy_es0_cnt <= (((hdmi_out0_driver_hdmi_phy_es0_cnt - $signed({1'd0, {(~hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es0_n0q_m}));
			end
		end
	end else begin
		hdmi_out0_driver_hdmi_phy_es0_out <= sync_f_array_muxed0;
		hdmi_out0_driver_hdmi_phy_es0_cnt <= 1'd0;
	end
	hdmi_out0_driver_hdmi_phy_es1_ce <= (~hdmi_out0_pix_rst);
	hdmi_out0_driver_hdmi_phy_es1_n1d <= (((((((hdmi_out0_driver_hdmi_phy_es1_d0[0] + hdmi_out0_driver_hdmi_phy_es1_d0[1]) + hdmi_out0_driver_hdmi_phy_es1_d0[2]) + hdmi_out0_driver_hdmi_phy_es1_d0[3]) + hdmi_out0_driver_hdmi_phy_es1_d0[4]) + hdmi_out0_driver_hdmi_phy_es1_d0[5]) + hdmi_out0_driver_hdmi_phy_es1_d0[6]) + hdmi_out0_driver_hdmi_phy_es1_d0[7]);
	hdmi_out0_driver_hdmi_phy_es1_d1 <= hdmi_out0_driver_hdmi_phy_es1_d0;
	hdmi_out0_driver_hdmi_phy_es1_q_m[0] <= hdmi_out0_driver_hdmi_phy_es1_d1[0];
	hdmi_out0_driver_hdmi_phy_es1_q_m[1] <= ((hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_q_m[2] <= ((((hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_q_m[3] <= ((((((hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_q_m[4] <= ((((((((hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_q_m[5] <= ((((((((((hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_q_m[6] <= ((((((((((((hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[6]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_q_m[7] <= ((((((((((((((hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[6]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es1_d1[7]) ^ hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_q_m[8] <= (~hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es1_n0q_m <= ((((((((~hdmi_out0_driver_hdmi_phy_es1_q_m[0]) + (~hdmi_out0_driver_hdmi_phy_es1_q_m[1])) + (~hdmi_out0_driver_hdmi_phy_es1_q_m[2])) + (~hdmi_out0_driver_hdmi_phy_es1_q_m[3])) + (~hdmi_out0_driver_hdmi_phy_es1_q_m[4])) + (~hdmi_out0_driver_hdmi_phy_es1_q_m[5])) + (~hdmi_out0_driver_hdmi_phy_es1_q_m[6])) + (~hdmi_out0_driver_hdmi_phy_es1_q_m[7]));
	hdmi_out0_driver_hdmi_phy_es1_n1q_m <= (((((((hdmi_out0_driver_hdmi_phy_es1_q_m[0] + hdmi_out0_driver_hdmi_phy_es1_q_m[1]) + hdmi_out0_driver_hdmi_phy_es1_q_m[2]) + hdmi_out0_driver_hdmi_phy_es1_q_m[3]) + hdmi_out0_driver_hdmi_phy_es1_q_m[4]) + hdmi_out0_driver_hdmi_phy_es1_q_m[5]) + hdmi_out0_driver_hdmi_phy_es1_q_m[6]) + hdmi_out0_driver_hdmi_phy_es1_q_m[7]);
	hdmi_out0_driver_hdmi_phy_es1_q_m_r <= hdmi_out0_driver_hdmi_phy_es1_q_m;
	hdmi_out0_driver_hdmi_phy_es1_new_c0 <= hdmi_out0_driver_hdmi_phy_es1_c;
	hdmi_out0_driver_hdmi_phy_es1_new_de0 <= hdmi_out0_driver_hdmi_phy_es1_de;
	hdmi_out0_driver_hdmi_phy_es1_new_c1 <= hdmi_out0_driver_hdmi_phy_es1_new_c0;
	hdmi_out0_driver_hdmi_phy_es1_new_de1 <= hdmi_out0_driver_hdmi_phy_es1_new_de0;
	hdmi_out0_driver_hdmi_phy_es1_new_c2 <= hdmi_out0_driver_hdmi_phy_es1_new_c1;
	hdmi_out0_driver_hdmi_phy_es1_new_de2 <= hdmi_out0_driver_hdmi_phy_es1_new_de1;
	if (hdmi_out0_driver_hdmi_phy_es1_new_de2) begin
		if (((hdmi_out0_driver_hdmi_phy_es1_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es1_n1q_m == hdmi_out0_driver_hdmi_phy_es1_n0q_m)}))) begin
			hdmi_out0_driver_hdmi_phy_es1_out[9] <= (~hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]);
			hdmi_out0_driver_hdmi_phy_es1_out[8] <= hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
			if (hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]) begin
				hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0];
				hdmi_out0_driver_hdmi_phy_es1_cnt <= ((hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n0q_m}));
			end else begin
				hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= (~hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0]);
				hdmi_out0_driver_hdmi_phy_es1_cnt <= ((hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n1q_m}));
			end
		end else begin
			if ((((~hdmi_out0_driver_hdmi_phy_es1_cnt[5]) & $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es1_n1q_m > hdmi_out0_driver_hdmi_phy_es1_n0q_m)})) | (hdmi_out0_driver_hdmi_phy_es1_cnt[5] & $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es1_n0q_m > hdmi_out0_driver_hdmi_phy_es1_n1q_m)})))) begin
				hdmi_out0_driver_hdmi_phy_es1_out[9] <= 1'd1;
				hdmi_out0_driver_hdmi_phy_es1_out[8] <= hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
				hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= (~hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0]);
				hdmi_out0_driver_hdmi_phy_es1_cnt <= (((hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, {hdmi_out0_driver_hdmi_phy_es1_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n1q_m}));
			end else begin
				hdmi_out0_driver_hdmi_phy_es1_out[9] <= 1'd0;
				hdmi_out0_driver_hdmi_phy_es1_out[8] <= hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
				hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0];
				hdmi_out0_driver_hdmi_phy_es1_cnt <= (((hdmi_out0_driver_hdmi_phy_es1_cnt - $signed({1'd0, {(~hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es1_n0q_m}));
			end
		end
	end else begin
		hdmi_out0_driver_hdmi_phy_es1_out <= sync_f_array_muxed1;
		hdmi_out0_driver_hdmi_phy_es1_cnt <= 1'd0;
	end
	hdmi_out0_driver_hdmi_phy_es2_ce <= (~hdmi_out0_pix_rst);
	hdmi_out0_driver_hdmi_phy_es2_n1d <= (((((((hdmi_out0_driver_hdmi_phy_es2_d0[0] + hdmi_out0_driver_hdmi_phy_es2_d0[1]) + hdmi_out0_driver_hdmi_phy_es2_d0[2]) + hdmi_out0_driver_hdmi_phy_es2_d0[3]) + hdmi_out0_driver_hdmi_phy_es2_d0[4]) + hdmi_out0_driver_hdmi_phy_es2_d0[5]) + hdmi_out0_driver_hdmi_phy_es2_d0[6]) + hdmi_out0_driver_hdmi_phy_es2_d0[7]);
	hdmi_out0_driver_hdmi_phy_es2_d1 <= hdmi_out0_driver_hdmi_phy_es2_d0;
	hdmi_out0_driver_hdmi_phy_es2_q_m[0] <= hdmi_out0_driver_hdmi_phy_es2_d1[0];
	hdmi_out0_driver_hdmi_phy_es2_q_m[1] <= ((hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_q_m[2] <= ((((hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_q_m[3] <= ((((((hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_q_m[4] <= ((((((((hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_q_m[5] <= ((((((((((hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_q_m[6] <= ((((((((((((hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[6]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_q_m[7] <= ((((((((((((((hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[6]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi_out0_driver_hdmi_phy_es2_d1[7]) ^ hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_q_m[8] <= (~hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi_out0_driver_hdmi_phy_es2_n0q_m <= ((((((((~hdmi_out0_driver_hdmi_phy_es2_q_m[0]) + (~hdmi_out0_driver_hdmi_phy_es2_q_m[1])) + (~hdmi_out0_driver_hdmi_phy_es2_q_m[2])) + (~hdmi_out0_driver_hdmi_phy_es2_q_m[3])) + (~hdmi_out0_driver_hdmi_phy_es2_q_m[4])) + (~hdmi_out0_driver_hdmi_phy_es2_q_m[5])) + (~hdmi_out0_driver_hdmi_phy_es2_q_m[6])) + (~hdmi_out0_driver_hdmi_phy_es2_q_m[7]));
	hdmi_out0_driver_hdmi_phy_es2_n1q_m <= (((((((hdmi_out0_driver_hdmi_phy_es2_q_m[0] + hdmi_out0_driver_hdmi_phy_es2_q_m[1]) + hdmi_out0_driver_hdmi_phy_es2_q_m[2]) + hdmi_out0_driver_hdmi_phy_es2_q_m[3]) + hdmi_out0_driver_hdmi_phy_es2_q_m[4]) + hdmi_out0_driver_hdmi_phy_es2_q_m[5]) + hdmi_out0_driver_hdmi_phy_es2_q_m[6]) + hdmi_out0_driver_hdmi_phy_es2_q_m[7]);
	hdmi_out0_driver_hdmi_phy_es2_q_m_r <= hdmi_out0_driver_hdmi_phy_es2_q_m;
	hdmi_out0_driver_hdmi_phy_es2_new_c0 <= hdmi_out0_driver_hdmi_phy_es2_c;
	hdmi_out0_driver_hdmi_phy_es2_new_de0 <= hdmi_out0_driver_hdmi_phy_es2_de;
	hdmi_out0_driver_hdmi_phy_es2_new_c1 <= hdmi_out0_driver_hdmi_phy_es2_new_c0;
	hdmi_out0_driver_hdmi_phy_es2_new_de1 <= hdmi_out0_driver_hdmi_phy_es2_new_de0;
	hdmi_out0_driver_hdmi_phy_es2_new_c2 <= hdmi_out0_driver_hdmi_phy_es2_new_c1;
	hdmi_out0_driver_hdmi_phy_es2_new_de2 <= hdmi_out0_driver_hdmi_phy_es2_new_de1;
	if (hdmi_out0_driver_hdmi_phy_es2_new_de2) begin
		if (((hdmi_out0_driver_hdmi_phy_es2_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es2_n1q_m == hdmi_out0_driver_hdmi_phy_es2_n0q_m)}))) begin
			hdmi_out0_driver_hdmi_phy_es2_out[9] <= (~hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]);
			hdmi_out0_driver_hdmi_phy_es2_out[8] <= hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
			if (hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]) begin
				hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0];
				hdmi_out0_driver_hdmi_phy_es2_cnt <= ((hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n0q_m}));
			end else begin
				hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= (~hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0]);
				hdmi_out0_driver_hdmi_phy_es2_cnt <= ((hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n1q_m}));
			end
		end else begin
			if ((((~hdmi_out0_driver_hdmi_phy_es2_cnt[5]) & $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es2_n1q_m > hdmi_out0_driver_hdmi_phy_es2_n0q_m)})) | (hdmi_out0_driver_hdmi_phy_es2_cnt[5] & $signed({1'd0, (hdmi_out0_driver_hdmi_phy_es2_n0q_m > hdmi_out0_driver_hdmi_phy_es2_n1q_m)})))) begin
				hdmi_out0_driver_hdmi_phy_es2_out[9] <= 1'd1;
				hdmi_out0_driver_hdmi_phy_es2_out[8] <= hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
				hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= (~hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0]);
				hdmi_out0_driver_hdmi_phy_es2_cnt <= (((hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, {hdmi_out0_driver_hdmi_phy_es2_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n1q_m}));
			end else begin
				hdmi_out0_driver_hdmi_phy_es2_out[9] <= 1'd0;
				hdmi_out0_driver_hdmi_phy_es2_out[8] <= hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
				hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0];
				hdmi_out0_driver_hdmi_phy_es2_cnt <= (((hdmi_out0_driver_hdmi_phy_es2_cnt - $signed({1'd0, {(~hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, hdmi_out0_driver_hdmi_phy_es2_n0q_m}));
			end
		end
	end else begin
		hdmi_out0_driver_hdmi_phy_es2_out <= sync_f_array_muxed2;
		hdmi_out0_driver_hdmi_phy_es2_cnt <= 1'd0;
	end
	if (hdmi_out0_pix_rst) begin
		hdmi_out0_dram_port_cmd_fifo_graycounter0_q <= 3'd0;
		hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary <= 3'd0;
		hdmi_out0_dram_port_rdata_fifo_graycounter1_q <= 5'd0;
		hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary <= 5'd0;
		hdmi_out0_dram_port_cmd_buffer_level <= 3'd0;
		hdmi_out0_dram_port_cmd_buffer_produce <= 2'd0;
		hdmi_out0_dram_port_cmd_buffer_consume <= 2'd0;
		hdmi_out0_dram_port_counter <= 3'd0;
		hdmi_out0_dram_port_rdata_buffer_valid_n <= 1'd0;
		hdmi_out0_dram_port_rdata_buffer_first_n <= 1'd0;
		hdmi_out0_dram_port_rdata_buffer_last_n <= 1'd0;
		hdmi_out0_dram_port_rdata_converter_converter_mux <= 3'd0;
		hdmi_out0_dram_port_rdata_chunk <= 8'd1;
		hdmi_out0_core_underflow_counter_status <= 32'd0;
		hdmi_out0_core_initiator_cdc_graycounter1_q <= 2'd0;
		hdmi_out0_core_initiator_cdc_graycounter1_q_binary <= 2'd0;
		hdmi_out0_core_timinggenerator_source_last <= 1'd0;
		hdmi_out0_core_timinggenerator_hactive <= 1'd0;
		hdmi_out0_core_timinggenerator_vactive <= 1'd0;
		hdmi_out0_core_timinggenerator_hcounter <= 12'd0;
		hdmi_out0_core_timinggenerator_vcounter <= 12'd0;
		hdmi_out0_core_dmareader_rsv_level <= 13'd0;
		hdmi_out0_core_dmareader_fifo_readable <= 1'd0;
		hdmi_out0_core_dmareader_fifo_level0 <= 13'd0;
		hdmi_out0_core_dmareader_fifo_produce <= 12'd0;
		hdmi_out0_core_dmareader_fifo_consume <= 12'd0;
		hdmi_out0_core_dmareader_offset <= 28'd0;
		hdmi_out0_core_underflow_counter <= 32'd0;
		hdmi_out0_driver_s7hdmioutclocking_ce <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es0_out <= 10'd0;
		hdmi_out0_driver_hdmi_phy_es0_d1 <= 8'd0;
		hdmi_out0_driver_hdmi_phy_es0_n1d <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es0_q_m <= 9'd0;
		hdmi_out0_driver_hdmi_phy_es0_q_m_r <= 9'd0;
		hdmi_out0_driver_hdmi_phy_es0_n0q_m <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es0_n1q_m <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es0_cnt <= 6'sd64;
		hdmi_out0_driver_hdmi_phy_es0_new_c0 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es0_new_de0 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es0_new_c1 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es0_new_de1 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es0_new_c2 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es0_new_de2 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es0_ce <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es1_out <= 10'd0;
		hdmi_out0_driver_hdmi_phy_es1_d1 <= 8'd0;
		hdmi_out0_driver_hdmi_phy_es1_n1d <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es1_q_m <= 9'd0;
		hdmi_out0_driver_hdmi_phy_es1_q_m_r <= 9'd0;
		hdmi_out0_driver_hdmi_phy_es1_n0q_m <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es1_n1q_m <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es1_cnt <= 6'sd64;
		hdmi_out0_driver_hdmi_phy_es1_new_c0 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es1_new_de0 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es1_new_c1 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es1_new_de1 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es1_new_c2 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es1_new_de2 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es1_ce <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es2_out <= 10'd0;
		hdmi_out0_driver_hdmi_phy_es2_d1 <= 8'd0;
		hdmi_out0_driver_hdmi_phy_es2_n1d <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es2_q_m <= 9'd0;
		hdmi_out0_driver_hdmi_phy_es2_q_m_r <= 9'd0;
		hdmi_out0_driver_hdmi_phy_es2_n0q_m <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es2_n1q_m <= 4'd0;
		hdmi_out0_driver_hdmi_phy_es2_cnt <= 6'sd64;
		hdmi_out0_driver_hdmi_phy_es2_new_c0 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es2_new_de0 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es2_new_c1 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es2_new_de1 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es2_new_c2 <= 2'd0;
		hdmi_out0_driver_hdmi_phy_es2_new_de2 <= 1'd0;
		hdmi_out0_driver_hdmi_phy_es2_ce <= 1'd0;
		hdmi_out0_resetinserter_y_fifo_level <= 3'd0;
		hdmi_out0_resetinserter_y_fifo_produce <= 2'd0;
		hdmi_out0_resetinserter_y_fifo_consume <= 2'd0;
		hdmi_out0_resetinserter_cb_fifo_level <= 3'd0;
		hdmi_out0_resetinserter_cb_fifo_produce <= 2'd0;
		hdmi_out0_resetinserter_cb_fifo_consume <= 2'd0;
		hdmi_out0_resetinserter_cr_fifo_level <= 3'd0;
		hdmi_out0_resetinserter_cr_fifo_produce <= 2'd0;
		hdmi_out0_resetinserter_cr_fifo_consume <= 2'd0;
		hdmi_out0_resetinserter_parity_in <= 1'd0;
		hdmi_out0_resetinserter_parity_out <= 1'd0;
		hdmi_out0_source_r <= 8'd0;
		hdmi_out0_source_g <= 8'd0;
		hdmi_out0_source_b <= 8'd0;
		hdmi_out0_record0_ycbcr_n_y <= 8'd0;
		hdmi_out0_record0_ycbcr_n_cb <= 8'd0;
		hdmi_out0_record0_ycbcr_n_cr <= 8'd0;
		hdmi_out0_record1_ycbcr_n_y <= 8'd0;
		hdmi_out0_record1_ycbcr_n_cb <= 8'd0;
		hdmi_out0_record1_ycbcr_n_cr <= 8'd0;
		hdmi_out0_record2_ycbcr_n_y <= 8'd0;
		hdmi_out0_record2_ycbcr_n_cb <= 8'd0;
		hdmi_out0_record2_ycbcr_n_cr <= 8'd0;
		hdmi_out0_record3_ycbcr_n_y <= 8'd0;
		hdmi_out0_record3_ycbcr_n_cb <= 8'd0;
		hdmi_out0_record3_ycbcr_n_cr <= 8'd0;
		hdmi_out0_cb_minus_coffset <= 9'sd512;
		hdmi_out0_cr_minus_coffset <= 9'sd512;
		hdmi_out0_y_minus_yoffset <= 9'sd512;
		hdmi_out0_cr_minus_coffset_mult_acoef <= 20'sd1048576;
		hdmi_out0_cb_minus_coffset_mult_bcoef <= 20'sd1048576;
		hdmi_out0_cr_minus_coffset_mult_ccoef <= 20'sd1048576;
		hdmi_out0_cb_minus_coffset_mult_dcoef <= 20'sd1048576;
		hdmi_out0_r <= 12'sd4096;
		hdmi_out0_g <= 12'sd4096;
		hdmi_out0_b <= 12'sd4096;
		hdmi_out0_valid_n0 <= 1'd0;
		hdmi_out0_valid_n1 <= 1'd0;
		hdmi_out0_valid_n2 <= 1'd0;
		hdmi_out0_valid_n3 <= 1'd0;
		hdmi_out0_first_n0 <= 1'd0;
		hdmi_out0_last_n0 <= 1'd0;
		hdmi_out0_first_n1 <= 1'd0;
		hdmi_out0_last_n1 <= 1'd0;
		hdmi_out0_first_n2 <= 1'd0;
		hdmi_out0_last_n2 <= 1'd0;
		hdmi_out0_first_n3 <= 1'd0;
		hdmi_out0_last_n3 <= 1'd0;
		hdmi_out0_next_s0 <= 1'd0;
		hdmi_out0_next_s1 <= 1'd0;
		hdmi_out0_next_s2 <= 1'd0;
		hdmi_out0_next_s3 <= 1'd0;
		hdmi_out0_next_s4 <= 1'd0;
		hdmi_out0_next_s5 <= 1'd0;
		hdmi_out0_next_s6 <= 1'd0;
		hdmi_out0_next_s7 <= 1'd0;
		hdmi_out0_next_s8 <= 1'd0;
		hdmi_out0_next_s9 <= 1'd0;
		hdmi_out0_next_s10 <= 1'd0;
		hdmi_out0_next_s11 <= 1'd0;
		hdmi_out0_next_s12 <= 1'd0;
		hdmi_out0_next_s13 <= 1'd0;
		hdmi_out0_next_s14 <= 1'd0;
		hdmi_out0_next_s15 <= 1'd0;
		hdmi_out0_next_s16 <= 1'd0;
		hdmi_out0_next_s17 <= 1'd0;
		hdmi_out0_de_r <= 1'd0;
		hdmi_out0_core_source_valid_d <= 1'd0;
		hdmi_out0_core_source_data_d <= 16'd0;
		videoout_state <= 1'd0;
	end
	xilinxmultiregimpl51_regs0 <= hdmi_out0_dram_port_cmd_fifo_graycounter1_q;
	xilinxmultiregimpl51_regs1 <= xilinxmultiregimpl51_regs0;
	xilinxmultiregimpl52_regs0 <= hdmi_out0_dram_port_rdata_fifo_graycounter0_q;
	xilinxmultiregimpl52_regs1 <= xilinxmultiregimpl52_regs0;
	xilinxmultiregimpl54_regs0 <= hdmi_out0_core_initiator_cdc_graycounter0_q;
	xilinxmultiregimpl54_regs1 <= xilinxmultiregimpl54_regs0;
	xilinxmultiregimpl57_regs0 <= hdmi_out0_core_toggle_i;
	xilinxmultiregimpl57_regs1 <= xilinxmultiregimpl57_regs0;
end

always @(posedge pix1p25x_clk) begin
	if (s7datacapture0_reset_lateness) begin
		s7datacapture0_lateness <= 8'd128;
	end else begin
		if (((~s7datacapture0_too_late) & (~s7datacapture0_too_early))) begin
			if (s7datacapture0_dec) begin
				s7datacapture0_lateness <= (s7datacapture0_lateness + 1'd1);
			end
			if (s7datacapture0_inc) begin
				s7datacapture0_lateness <= (s7datacapture0_lateness - 1'd1);
			end
		end
	end
	s7datacapture0_mdata_d <= s7datacapture0_mdata;
	s7datacapture0_do_delay_rst_toggle_o_r <= s7datacapture0_do_delay_rst_toggle_o;
	s7datacapture0_do_delay_master_inc_toggle_o_r <= s7datacapture0_do_delay_master_inc_toggle_o;
	s7datacapture0_do_delay_master_dec_toggle_o_r <= s7datacapture0_do_delay_master_dec_toggle_o;
	s7datacapture0_do_delay_slave_inc_toggle_o_r <= s7datacapture0_do_delay_slave_inc_toggle_o;
	s7datacapture0_do_delay_slave_dec_toggle_o_r <= s7datacapture0_do_delay_slave_dec_toggle_o;
	s7datacapture0_do_reset_lateness_toggle_o_r <= s7datacapture0_do_reset_lateness_toggle_o;
	if (s7datacapture1_reset_lateness) begin
		s7datacapture1_lateness <= 8'd128;
	end else begin
		if (((~s7datacapture1_too_late) & (~s7datacapture1_too_early))) begin
			if (s7datacapture1_dec) begin
				s7datacapture1_lateness <= (s7datacapture1_lateness + 1'd1);
			end
			if (s7datacapture1_inc) begin
				s7datacapture1_lateness <= (s7datacapture1_lateness - 1'd1);
			end
		end
	end
	s7datacapture1_mdata_d <= s7datacapture1_mdata;
	s7datacapture1_do_delay_rst_toggle_o_r <= s7datacapture1_do_delay_rst_toggle_o;
	s7datacapture1_do_delay_master_inc_toggle_o_r <= s7datacapture1_do_delay_master_inc_toggle_o;
	s7datacapture1_do_delay_master_dec_toggle_o_r <= s7datacapture1_do_delay_master_dec_toggle_o;
	s7datacapture1_do_delay_slave_inc_toggle_o_r <= s7datacapture1_do_delay_slave_inc_toggle_o;
	s7datacapture1_do_delay_slave_dec_toggle_o_r <= s7datacapture1_do_delay_slave_dec_toggle_o;
	s7datacapture1_do_reset_lateness_toggle_o_r <= s7datacapture1_do_reset_lateness_toggle_o;
	if (s7datacapture2_reset_lateness) begin
		s7datacapture2_lateness <= 8'd128;
	end else begin
		if (((~s7datacapture2_too_late) & (~s7datacapture2_too_early))) begin
			if (s7datacapture2_dec) begin
				s7datacapture2_lateness <= (s7datacapture2_lateness + 1'd1);
			end
			if (s7datacapture2_inc) begin
				s7datacapture2_lateness <= (s7datacapture2_lateness - 1'd1);
			end
		end
	end
	s7datacapture2_mdata_d <= s7datacapture2_mdata;
	s7datacapture2_do_delay_rst_toggle_o_r <= s7datacapture2_do_delay_rst_toggle_o;
	s7datacapture2_do_delay_master_inc_toggle_o_r <= s7datacapture2_do_delay_master_inc_toggle_o;
	s7datacapture2_do_delay_master_dec_toggle_o_r <= s7datacapture2_do_delay_master_dec_toggle_o;
	s7datacapture2_do_delay_slave_inc_toggle_o_r <= s7datacapture2_do_delay_slave_inc_toggle_o;
	s7datacapture2_do_delay_slave_dec_toggle_o_r <= s7datacapture2_do_delay_slave_dec_toggle_o;
	s7datacapture2_do_reset_lateness_toggle_o_r <= s7datacapture2_do_reset_lateness_toggle_o;
	if (pix1p25x_rst) begin
		s7datacapture0_mdata_d <= 8'd0;
		s7datacapture0_lateness <= 8'd128;
		s7datacapture1_mdata_d <= 8'd0;
		s7datacapture1_lateness <= 8'd128;
		s7datacapture2_mdata_d <= 8'd0;
		s7datacapture2_lateness <= 8'd128;
	end
	xilinxmultiregimpl11_regs0 <= s7datacapture0_do_delay_rst_toggle_i;
	xilinxmultiregimpl11_regs1 <= xilinxmultiregimpl11_regs0;
	xilinxmultiregimpl12_regs0 <= s7datacapture0_do_delay_master_inc_toggle_i;
	xilinxmultiregimpl12_regs1 <= xilinxmultiregimpl12_regs0;
	xilinxmultiregimpl13_regs0 <= s7datacapture0_do_delay_master_dec_toggle_i;
	xilinxmultiregimpl13_regs1 <= xilinxmultiregimpl13_regs0;
	xilinxmultiregimpl14_regs0 <= s7datacapture0_do_delay_slave_inc_toggle_i;
	xilinxmultiregimpl14_regs1 <= xilinxmultiregimpl14_regs0;
	xilinxmultiregimpl15_regs0 <= s7datacapture0_do_delay_slave_dec_toggle_i;
	xilinxmultiregimpl15_regs1 <= xilinxmultiregimpl15_regs0;
	xilinxmultiregimpl17_regs0 <= s7datacapture0_do_reset_lateness_toggle_i;
	xilinxmultiregimpl17_regs1 <= xilinxmultiregimpl17_regs0;
	xilinxmultiregimpl21_regs0 <= s7datacapture1_do_delay_rst_toggle_i;
	xilinxmultiregimpl21_regs1 <= xilinxmultiregimpl21_regs0;
	xilinxmultiregimpl22_regs0 <= s7datacapture1_do_delay_master_inc_toggle_i;
	xilinxmultiregimpl22_regs1 <= xilinxmultiregimpl22_regs0;
	xilinxmultiregimpl23_regs0 <= s7datacapture1_do_delay_master_dec_toggle_i;
	xilinxmultiregimpl23_regs1 <= xilinxmultiregimpl23_regs0;
	xilinxmultiregimpl24_regs0 <= s7datacapture1_do_delay_slave_inc_toggle_i;
	xilinxmultiregimpl24_regs1 <= xilinxmultiregimpl24_regs0;
	xilinxmultiregimpl25_regs0 <= s7datacapture1_do_delay_slave_dec_toggle_i;
	xilinxmultiregimpl25_regs1 <= xilinxmultiregimpl25_regs0;
	xilinxmultiregimpl27_regs0 <= s7datacapture1_do_reset_lateness_toggle_i;
	xilinxmultiregimpl27_regs1 <= xilinxmultiregimpl27_regs0;
	xilinxmultiregimpl31_regs0 <= s7datacapture2_do_delay_rst_toggle_i;
	xilinxmultiregimpl31_regs1 <= xilinxmultiregimpl31_regs0;
	xilinxmultiregimpl32_regs0 <= s7datacapture2_do_delay_master_inc_toggle_i;
	xilinxmultiregimpl32_regs1 <= xilinxmultiregimpl32_regs0;
	xilinxmultiregimpl33_regs0 <= s7datacapture2_do_delay_master_dec_toggle_i;
	xilinxmultiregimpl33_regs1 <= xilinxmultiregimpl33_regs0;
	xilinxmultiregimpl34_regs0 <= s7datacapture2_do_delay_slave_inc_toggle_i;
	xilinxmultiregimpl34_regs1 <= xilinxmultiregimpl34_regs0;
	xilinxmultiregimpl35_regs0 <= s7datacapture2_do_delay_slave_dec_toggle_i;
	xilinxmultiregimpl35_regs1 <= xilinxmultiregimpl35_regs0;
	xilinxmultiregimpl37_regs0 <= s7datacapture2_do_reset_lateness_toggle_i;
	xilinxmultiregimpl37_regs1 <= xilinxmultiregimpl37_regs0;
end

always @(posedge sys_clk) begin
	videosoc_videosoc_rom_bus_ack <= 1'd0;
	if (((videosoc_videosoc_rom_bus_cyc & videosoc_videosoc_rom_bus_stb) & (~videosoc_videosoc_rom_bus_ack))) begin
		videosoc_videosoc_rom_bus_ack <= 1'd1;
	end
	videosoc_videosoc_sram_bus_ack <= 1'd0;
	if (((videosoc_videosoc_sram_bus_cyc & videosoc_videosoc_sram_bus_stb) & (~videosoc_videosoc_sram_bus_ack))) begin
		videosoc_videosoc_sram_bus_ack <= 1'd1;
	end
	videosoc_videosoc_interface_we <= 1'd0;
	videosoc_videosoc_interface_dat_w <= videosoc_videosoc_bus_wishbone_dat_w;
	videosoc_videosoc_interface_adr <= videosoc_videosoc_bus_wishbone_adr;
	videosoc_videosoc_bus_wishbone_dat_r <= videosoc_videosoc_interface_dat_r;
	if ((videosoc_videosoc_counter == 1'd1)) begin
		videosoc_videosoc_interface_we <= videosoc_videosoc_bus_wishbone_we;
	end
	if ((videosoc_videosoc_counter == 2'd2)) begin
		videosoc_videosoc_bus_wishbone_ack <= 1'd1;
	end
	if ((videosoc_videosoc_counter == 2'd3)) begin
		videosoc_videosoc_bus_wishbone_ack <= 1'd0;
	end
	if ((videosoc_videosoc_counter != 1'd0)) begin
		videosoc_videosoc_counter <= (videosoc_videosoc_counter + 1'd1);
	end else begin
		if ((videosoc_videosoc_bus_wishbone_cyc & videosoc_videosoc_bus_wishbone_stb)) begin
			videosoc_videosoc_counter <= 1'd1;
		end
	end
	if (videosoc_videosoc_en_storage) begin
		if ((videosoc_videosoc_value == 1'd0)) begin
			videosoc_videosoc_value <= videosoc_videosoc_reload_storage;
		end else begin
			videosoc_videosoc_value <= (videosoc_videosoc_value - 1'd1);
		end
	end else begin
		videosoc_videosoc_value <= videosoc_videosoc_load_storage;
	end
	if (videosoc_videosoc_update_value_re) begin
		videosoc_videosoc_value_status <= videosoc_videosoc_value;
	end
	if (videosoc_videosoc_zero_clear) begin
		videosoc_videosoc_zero_pending <= 1'd0;
	end
	videosoc_videosoc_zero_old_trigger <= videosoc_videosoc_zero_trigger;
	if (((~videosoc_videosoc_zero_trigger) & videosoc_videosoc_zero_old_trigger)) begin
		videosoc_videosoc_zero_pending <= 1'd1;
	end
	if (videosoc_uart_tx_clear) begin
		videosoc_uart_tx_pending <= 1'd0;
	end
	videosoc_uart_tx_old_trigger <= videosoc_uart_tx_trigger;
	if (((~videosoc_uart_tx_trigger) & videosoc_uart_tx_old_trigger)) begin
		videosoc_uart_tx_pending <= 1'd1;
	end
	if (videosoc_uart_rx_clear) begin
		videosoc_uart_rx_pending <= 1'd0;
	end
	videosoc_uart_rx_old_trigger <= videosoc_uart_rx_trigger;
	if (((~videosoc_uart_rx_trigger) & videosoc_uart_rx_old_trigger)) begin
		videosoc_uart_rx_pending <= 1'd1;
	end
	if (((videosoc_uart_tx_fifo_syncfifo_we & videosoc_uart_tx_fifo_syncfifo_writable) & (~videosoc_uart_tx_fifo_replace))) begin
		videosoc_uart_tx_fifo_produce <= (videosoc_uart_tx_fifo_produce + 1'd1);
	end
	if (videosoc_uart_tx_fifo_do_read) begin
		videosoc_uart_tx_fifo_consume <= (videosoc_uart_tx_fifo_consume + 1'd1);
	end
	if (((videosoc_uart_tx_fifo_syncfifo_we & videosoc_uart_tx_fifo_syncfifo_writable) & (~videosoc_uart_tx_fifo_replace))) begin
		if ((~videosoc_uart_tx_fifo_do_read)) begin
			videosoc_uart_tx_fifo_level <= (videosoc_uart_tx_fifo_level + 1'd1);
		end
	end else begin
		if (videosoc_uart_tx_fifo_do_read) begin
			videosoc_uart_tx_fifo_level <= (videosoc_uart_tx_fifo_level - 1'd1);
		end
	end
	if (((videosoc_uart_rx_fifo_syncfifo_we & videosoc_uart_rx_fifo_syncfifo_writable) & (~videosoc_uart_rx_fifo_replace))) begin
		videosoc_uart_rx_fifo_produce <= (videosoc_uart_rx_fifo_produce + 1'd1);
	end
	if (videosoc_uart_rx_fifo_do_read) begin
		videosoc_uart_rx_fifo_consume <= (videosoc_uart_rx_fifo_consume + 1'd1);
	end
	if (((videosoc_uart_rx_fifo_syncfifo_we & videosoc_uart_rx_fifo_syncfifo_writable) & (~videosoc_uart_rx_fifo_replace))) begin
		if ((~videosoc_uart_rx_fifo_do_read)) begin
			videosoc_uart_rx_fifo_level <= (videosoc_uart_rx_fifo_level + 1'd1);
		end
	end else begin
		if (videosoc_uart_rx_fifo_do_read) begin
			videosoc_uart_rx_fifo_level <= (videosoc_uart_rx_fifo_level - 1'd1);
		end
	end
	if (videosoc_bridge_byte_counter_reset) begin
		videosoc_bridge_byte_counter <= 1'd0;
	end else begin
		if (videosoc_bridge_byte_counter_ce) begin
			videosoc_bridge_byte_counter <= (videosoc_bridge_byte_counter + 1'd1);
		end
	end
	if (videosoc_bridge_word_counter_reset) begin
		videosoc_bridge_word_counter <= 1'd0;
	end else begin
		if (videosoc_bridge_word_counter_ce) begin
			videosoc_bridge_word_counter <= (videosoc_bridge_word_counter + 1'd1);
		end
	end
	if (videosoc_bridge_cmd_ce) begin
		videosoc_bridge_cmd <= videosoc_rs232phyinterface1_source_payload_data;
	end
	if (videosoc_bridge_length_ce) begin
		videosoc_bridge_length <= videosoc_rs232phyinterface1_source_payload_data;
	end
	if (videosoc_bridge_address_ce) begin
		videosoc_bridge_address <= {videosoc_bridge_address[23:0], videosoc_rs232phyinterface1_source_payload_data};
	end
	if (videosoc_bridge_rx_data_ce) begin
		videosoc_bridge_data <= {videosoc_bridge_data[23:0], videosoc_rs232phyinterface1_source_payload_data};
	end else begin
		if (videosoc_bridge_tx_data_ce) begin
			videosoc_bridge_data <= videosoc_bridge_wishbone_dat_r;
		end
	end
	wishbonestreamingbridge_state <= wishbonestreamingbridge_next_state;
	if (videosoc_bridge_reset) begin
		wishbonestreamingbridge_state <= 3'd0;
	end
	if (videosoc_bridge_wait) begin
		if ((~videosoc_bridge_done)) begin
			videosoc_bridge_count <= (videosoc_bridge_count - 1'd1);
		end
	end else begin
		videosoc_bridge_count <= 24'd10000000;
	end
	videosoc_uart_phy_sink_ready <= 1'd0;
	if (((videosoc_uart_phy_sink_valid & (~videosoc_uart_phy_tx_busy)) & (~videosoc_uart_phy_sink_ready))) begin
		videosoc_uart_phy_tx_reg <= videosoc_uart_phy_sink_payload_data;
		videosoc_uart_phy_tx_bitcount <= 1'd0;
		videosoc_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((videosoc_uart_phy_uart_clk_txen & videosoc_uart_phy_tx_busy)) begin
			videosoc_uart_phy_tx_bitcount <= (videosoc_uart_phy_tx_bitcount + 1'd1);
			if ((videosoc_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((videosoc_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					videosoc_uart_phy_tx_busy <= 1'd0;
					videosoc_uart_phy_sink_ready <= 1'd1;
				end else begin
					serial_tx <= videosoc_uart_phy_tx_reg[0];
					videosoc_uart_phy_tx_reg <= {1'd0, videosoc_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (videosoc_uart_phy_tx_busy) begin
		{videosoc_uart_phy_uart_clk_txen, videosoc_uart_phy_phase_accumulator_tx} <= (videosoc_uart_phy_phase_accumulator_tx + videosoc_uart_phy_storage);
	end else begin
		{videosoc_uart_phy_uart_clk_txen, videosoc_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	videosoc_uart_phy_source_valid <= 1'd0;
	videosoc_uart_phy_rx_r <= videosoc_uart_phy_rx;
	if ((~videosoc_uart_phy_rx_busy)) begin
		if (((~videosoc_uart_phy_rx) & videosoc_uart_phy_rx_r)) begin
			videosoc_uart_phy_rx_busy <= 1'd1;
			videosoc_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (videosoc_uart_phy_uart_clk_rxen) begin
			videosoc_uart_phy_rx_bitcount <= (videosoc_uart_phy_rx_bitcount + 1'd1);
			if ((videosoc_uart_phy_rx_bitcount == 1'd0)) begin
				if (videosoc_uart_phy_rx) begin
					videosoc_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((videosoc_uart_phy_rx_bitcount == 4'd9)) begin
					videosoc_uart_phy_rx_busy <= 1'd0;
					if (videosoc_uart_phy_rx) begin
						videosoc_uart_phy_source_payload_data <= videosoc_uart_phy_rx_reg;
						videosoc_uart_phy_source_valid <= 1'd1;
					end
				end else begin
					videosoc_uart_phy_rx_reg <= {videosoc_uart_phy_rx, videosoc_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (videosoc_uart_phy_rx_busy) begin
		{videosoc_uart_phy_uart_clk_rxen, videosoc_uart_phy_phase_accumulator_rx} <= (videosoc_uart_phy_phase_accumulator_rx + videosoc_uart_phy_storage);
	end else begin
		{videosoc_uart_phy_uart_clk_rxen, videosoc_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if ((videosoc_info_dna_cnt < 7'd114)) begin
		videosoc_info_dna_cnt <= (videosoc_info_dna_cnt + 1'd1);
		if (videosoc_info_dna_cnt[0]) begin
			videosoc_info_dna_status <= {videosoc_info_dna_status, videosoc_info_dna_do};
		end
	end
	if (videosoc_info_drdy) begin
		case (videosoc_info_channel)
			1'd0: begin
				videosoc_info_temperature_status <= (videosoc_info_data >>> 3'd4);
			end
			1'd1: begin
				videosoc_info_vccint_status <= (videosoc_info_data >>> 3'd4);
			end
			2'd2: begin
				videosoc_info_vccaux_status <= (videosoc_info_data >>> 3'd4);
			end
			3'd6: begin
				videosoc_info_vccbram_status <= (videosoc_info_data >>> 3'd4);
			end
		endcase
	end
	if (videosoc_oled_spimaster_set_clk) begin
		videosoc_oled_spi_pads_clk <= videosoc_oled_spimaster_enable_cs;
	end
	if (videosoc_oled_spimaster_clr_clk) begin
		videosoc_oled_spi_pads_clk <= 1'd0;
		videosoc_oled_spimaster_i <= 1'd0;
	end else begin
		videosoc_oled_spimaster_i <= (videosoc_oled_spimaster_i + 1'd1);
	end
	if (videosoc_oled_spimaster_clr_cnt) begin
		videosoc_oled_spimaster_cnt <= 1'd0;
	end else begin
		if (videosoc_oled_spimaster_inc_cnt) begin
			videosoc_oled_spimaster_cnt <= (videosoc_oled_spimaster_cnt + 1'd1);
		end
	end
	if (videosoc_oled_spimaster_start) begin
		videosoc_oled_spimaster_sr_mosi <= videosoc_oled_spimaster_mosi_storage;
	end else begin
		if ((videosoc_oled_spimaster_set_clk & videosoc_oled_spimaster_enable_shift)) begin
			videosoc_oled_spimaster_sr_mosi <= {videosoc_oled_spimaster_sr_mosi[6:0], videosoc_oled_spimaster};
		end else begin
			if (videosoc_oled_spimaster_clr_clk) begin
				videosoc_oled_spi_pads_mosi <= videosoc_oled_spimaster_sr_mosi[7];
			end
		end
	end
	oled_state <= oled_next_state;
	videosoc_ddrphy_n_rddata_en0 <= videosoc_ddrphy_dfi_p0_rddata_en;
	videosoc_ddrphy_n_rddata_en1 <= videosoc_ddrphy_n_rddata_en0;
	videosoc_ddrphy_n_rddata_en2 <= videosoc_ddrphy_n_rddata_en1;
	videosoc_ddrphy_n_rddata_en3 <= videosoc_ddrphy_n_rddata_en2;
	videosoc_ddrphy_n_rddata_en4 <= videosoc_ddrphy_n_rddata_en3;
	videosoc_ddrphy_dfi_p0_rddata_valid <= videosoc_ddrphy_n_rddata_en4;
	videosoc_ddrphy_dfi_p1_rddata_valid <= videosoc_ddrphy_n_rddata_en4;
	videosoc_ddrphy_dfi_p2_rddata_valid <= videosoc_ddrphy_n_rddata_en4;
	videosoc_ddrphy_dfi_p3_rddata_valid <= videosoc_ddrphy_n_rddata_en4;
	videosoc_ddrphy_last_wrdata_en <= {videosoc_ddrphy_last_wrdata_en[2:0], videosoc_ddrphy_dfi_p2_wrdata_en};
	videosoc_ddrphy_oe_dqs <= videosoc_ddrphy_oe;
	videosoc_ddrphy_oe_dq <= videosoc_ddrphy_oe;
	if (videosoc_sdram_inti_p0_rddata_valid) begin
		videosoc_sdram_phaseinjector0_status <= videosoc_sdram_inti_p0_rddata;
	end
	if (videosoc_sdram_inti_p1_rddata_valid) begin
		videosoc_sdram_phaseinjector1_status <= videosoc_sdram_inti_p1_rddata;
	end
	if (videosoc_sdram_inti_p2_rddata_valid) begin
		videosoc_sdram_phaseinjector2_status <= videosoc_sdram_inti_p2_rddata;
	end
	if (videosoc_sdram_inti_p3_rddata_valid) begin
		videosoc_sdram_phaseinjector3_status <= videosoc_sdram_inti_p3_rddata;
	end
	videosoc_sdram_cmd_payload_a <= 11'd1024;
	videosoc_sdram_cmd_payload_ba <= 1'd0;
	videosoc_sdram_cmd_payload_cas <= 1'd0;
	videosoc_sdram_cmd_payload_ras <= 1'd0;
	videosoc_sdram_cmd_payload_we <= 1'd0;
	videosoc_sdram_seq_done <= 1'd0;
	if ((videosoc_sdram_counter == 1'd1)) begin
		videosoc_sdram_cmd_payload_ras <= 1'd1;
		videosoc_sdram_cmd_payload_we <= 1'd1;
	end
	if ((videosoc_sdram_counter == 3'd4)) begin
		videosoc_sdram_cmd_payload_cas <= 1'd1;
		videosoc_sdram_cmd_payload_ras <= 1'd1;
	end
	if ((videosoc_sdram_counter == 5'd31)) begin
		videosoc_sdram_seq_done <= 1'd1;
	end
	if ((videosoc_sdram_counter != 1'd0)) begin
		videosoc_sdram_counter <= (videosoc_sdram_counter + 1'd1);
	end else begin
		if (videosoc_sdram_seq_start) begin
			videosoc_sdram_counter <= 1'd1;
		end
	end
	if (videosoc_sdram_wait) begin
		if ((~videosoc_sdram_done)) begin
			videosoc_sdram_count <= (videosoc_sdram_count - 1'd1);
		end
	end else begin
		videosoc_sdram_count <= 10'd782;
	end
	refresher_state <= refresher_next_state;
	if (videosoc_sdram_bankmachine0_track_close) begin
		videosoc_sdram_bankmachine0_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine0_track_open) begin
			videosoc_sdram_bankmachine0_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine0_openrow <= videosoc_sdram_bankmachine0_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine0_syncfifo0_we & videosoc_sdram_bankmachine0_syncfifo0_writable) & (~videosoc_sdram_bankmachine0_replace))) begin
		videosoc_sdram_bankmachine0_produce <= (videosoc_sdram_bankmachine0_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine0_do_read) begin
		videosoc_sdram_bankmachine0_consume <= (videosoc_sdram_bankmachine0_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine0_syncfifo0_we & videosoc_sdram_bankmachine0_syncfifo0_writable) & (~videosoc_sdram_bankmachine0_replace))) begin
		if ((~videosoc_sdram_bankmachine0_do_read)) begin
			videosoc_sdram_bankmachine0_level <= (videosoc_sdram_bankmachine0_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine0_do_read) begin
			videosoc_sdram_bankmachine0_level <= (videosoc_sdram_bankmachine0_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine0_wait) begin
		if ((~videosoc_sdram_bankmachine0_done)) begin
			videosoc_sdram_bankmachine0_count <= (videosoc_sdram_bankmachine0_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine0_count <= 3'd5;
	end
	bankmachine0_state <= bankmachine0_next_state;
	if (videosoc_sdram_bankmachine1_track_close) begin
		videosoc_sdram_bankmachine1_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine1_track_open) begin
			videosoc_sdram_bankmachine1_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine1_openrow <= videosoc_sdram_bankmachine1_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine1_syncfifo1_we & videosoc_sdram_bankmachine1_syncfifo1_writable) & (~videosoc_sdram_bankmachine1_replace))) begin
		videosoc_sdram_bankmachine1_produce <= (videosoc_sdram_bankmachine1_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine1_do_read) begin
		videosoc_sdram_bankmachine1_consume <= (videosoc_sdram_bankmachine1_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine1_syncfifo1_we & videosoc_sdram_bankmachine1_syncfifo1_writable) & (~videosoc_sdram_bankmachine1_replace))) begin
		if ((~videosoc_sdram_bankmachine1_do_read)) begin
			videosoc_sdram_bankmachine1_level <= (videosoc_sdram_bankmachine1_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine1_do_read) begin
			videosoc_sdram_bankmachine1_level <= (videosoc_sdram_bankmachine1_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine1_wait) begin
		if ((~videosoc_sdram_bankmachine1_done)) begin
			videosoc_sdram_bankmachine1_count <= (videosoc_sdram_bankmachine1_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine1_count <= 3'd5;
	end
	bankmachine1_state <= bankmachine1_next_state;
	if (videosoc_sdram_bankmachine2_track_close) begin
		videosoc_sdram_bankmachine2_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine2_track_open) begin
			videosoc_sdram_bankmachine2_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine2_openrow <= videosoc_sdram_bankmachine2_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine2_syncfifo2_we & videosoc_sdram_bankmachine2_syncfifo2_writable) & (~videosoc_sdram_bankmachine2_replace))) begin
		videosoc_sdram_bankmachine2_produce <= (videosoc_sdram_bankmachine2_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine2_do_read) begin
		videosoc_sdram_bankmachine2_consume <= (videosoc_sdram_bankmachine2_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine2_syncfifo2_we & videosoc_sdram_bankmachine2_syncfifo2_writable) & (~videosoc_sdram_bankmachine2_replace))) begin
		if ((~videosoc_sdram_bankmachine2_do_read)) begin
			videosoc_sdram_bankmachine2_level <= (videosoc_sdram_bankmachine2_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine2_do_read) begin
			videosoc_sdram_bankmachine2_level <= (videosoc_sdram_bankmachine2_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine2_wait) begin
		if ((~videosoc_sdram_bankmachine2_done)) begin
			videosoc_sdram_bankmachine2_count <= (videosoc_sdram_bankmachine2_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine2_count <= 3'd5;
	end
	bankmachine2_state <= bankmachine2_next_state;
	if (videosoc_sdram_bankmachine3_track_close) begin
		videosoc_sdram_bankmachine3_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine3_track_open) begin
			videosoc_sdram_bankmachine3_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine3_openrow <= videosoc_sdram_bankmachine3_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine3_syncfifo3_we & videosoc_sdram_bankmachine3_syncfifo3_writable) & (~videosoc_sdram_bankmachine3_replace))) begin
		videosoc_sdram_bankmachine3_produce <= (videosoc_sdram_bankmachine3_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine3_do_read) begin
		videosoc_sdram_bankmachine3_consume <= (videosoc_sdram_bankmachine3_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine3_syncfifo3_we & videosoc_sdram_bankmachine3_syncfifo3_writable) & (~videosoc_sdram_bankmachine3_replace))) begin
		if ((~videosoc_sdram_bankmachine3_do_read)) begin
			videosoc_sdram_bankmachine3_level <= (videosoc_sdram_bankmachine3_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine3_do_read) begin
			videosoc_sdram_bankmachine3_level <= (videosoc_sdram_bankmachine3_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine3_wait) begin
		if ((~videosoc_sdram_bankmachine3_done)) begin
			videosoc_sdram_bankmachine3_count <= (videosoc_sdram_bankmachine3_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine3_count <= 3'd5;
	end
	bankmachine3_state <= bankmachine3_next_state;
	if (videosoc_sdram_bankmachine4_track_close) begin
		videosoc_sdram_bankmachine4_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine4_track_open) begin
			videosoc_sdram_bankmachine4_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine4_openrow <= videosoc_sdram_bankmachine4_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine4_syncfifo4_we & videosoc_sdram_bankmachine4_syncfifo4_writable) & (~videosoc_sdram_bankmachine4_replace))) begin
		videosoc_sdram_bankmachine4_produce <= (videosoc_sdram_bankmachine4_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine4_do_read) begin
		videosoc_sdram_bankmachine4_consume <= (videosoc_sdram_bankmachine4_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine4_syncfifo4_we & videosoc_sdram_bankmachine4_syncfifo4_writable) & (~videosoc_sdram_bankmachine4_replace))) begin
		if ((~videosoc_sdram_bankmachine4_do_read)) begin
			videosoc_sdram_bankmachine4_level <= (videosoc_sdram_bankmachine4_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine4_do_read) begin
			videosoc_sdram_bankmachine4_level <= (videosoc_sdram_bankmachine4_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine4_wait) begin
		if ((~videosoc_sdram_bankmachine4_done)) begin
			videosoc_sdram_bankmachine4_count <= (videosoc_sdram_bankmachine4_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine4_count <= 3'd5;
	end
	bankmachine4_state <= bankmachine4_next_state;
	if (videosoc_sdram_bankmachine5_track_close) begin
		videosoc_sdram_bankmachine5_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine5_track_open) begin
			videosoc_sdram_bankmachine5_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine5_openrow <= videosoc_sdram_bankmachine5_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine5_syncfifo5_we & videosoc_sdram_bankmachine5_syncfifo5_writable) & (~videosoc_sdram_bankmachine5_replace))) begin
		videosoc_sdram_bankmachine5_produce <= (videosoc_sdram_bankmachine5_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine5_do_read) begin
		videosoc_sdram_bankmachine5_consume <= (videosoc_sdram_bankmachine5_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine5_syncfifo5_we & videosoc_sdram_bankmachine5_syncfifo5_writable) & (~videosoc_sdram_bankmachine5_replace))) begin
		if ((~videosoc_sdram_bankmachine5_do_read)) begin
			videosoc_sdram_bankmachine5_level <= (videosoc_sdram_bankmachine5_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine5_do_read) begin
			videosoc_sdram_bankmachine5_level <= (videosoc_sdram_bankmachine5_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine5_wait) begin
		if ((~videosoc_sdram_bankmachine5_done)) begin
			videosoc_sdram_bankmachine5_count <= (videosoc_sdram_bankmachine5_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine5_count <= 3'd5;
	end
	bankmachine5_state <= bankmachine5_next_state;
	if (videosoc_sdram_bankmachine6_track_close) begin
		videosoc_sdram_bankmachine6_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine6_track_open) begin
			videosoc_sdram_bankmachine6_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine6_openrow <= videosoc_sdram_bankmachine6_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine6_syncfifo6_we & videosoc_sdram_bankmachine6_syncfifo6_writable) & (~videosoc_sdram_bankmachine6_replace))) begin
		videosoc_sdram_bankmachine6_produce <= (videosoc_sdram_bankmachine6_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine6_do_read) begin
		videosoc_sdram_bankmachine6_consume <= (videosoc_sdram_bankmachine6_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine6_syncfifo6_we & videosoc_sdram_bankmachine6_syncfifo6_writable) & (~videosoc_sdram_bankmachine6_replace))) begin
		if ((~videosoc_sdram_bankmachine6_do_read)) begin
			videosoc_sdram_bankmachine6_level <= (videosoc_sdram_bankmachine6_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine6_do_read) begin
			videosoc_sdram_bankmachine6_level <= (videosoc_sdram_bankmachine6_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine6_wait) begin
		if ((~videosoc_sdram_bankmachine6_done)) begin
			videosoc_sdram_bankmachine6_count <= (videosoc_sdram_bankmachine6_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine6_count <= 3'd5;
	end
	bankmachine6_state <= bankmachine6_next_state;
	if (videosoc_sdram_bankmachine7_track_close) begin
		videosoc_sdram_bankmachine7_has_openrow <= 1'd0;
	end else begin
		if (videosoc_sdram_bankmachine7_track_open) begin
			videosoc_sdram_bankmachine7_has_openrow <= 1'd1;
			videosoc_sdram_bankmachine7_openrow <= videosoc_sdram_bankmachine7_source_payload_adr[21:7];
		end
	end
	if (((videosoc_sdram_bankmachine7_syncfifo7_we & videosoc_sdram_bankmachine7_syncfifo7_writable) & (~videosoc_sdram_bankmachine7_replace))) begin
		videosoc_sdram_bankmachine7_produce <= (videosoc_sdram_bankmachine7_produce + 1'd1);
	end
	if (videosoc_sdram_bankmachine7_do_read) begin
		videosoc_sdram_bankmachine7_consume <= (videosoc_sdram_bankmachine7_consume + 1'd1);
	end
	if (((videosoc_sdram_bankmachine7_syncfifo7_we & videosoc_sdram_bankmachine7_syncfifo7_writable) & (~videosoc_sdram_bankmachine7_replace))) begin
		if ((~videosoc_sdram_bankmachine7_do_read)) begin
			videosoc_sdram_bankmachine7_level <= (videosoc_sdram_bankmachine7_level + 1'd1);
		end
	end else begin
		if (videosoc_sdram_bankmachine7_do_read) begin
			videosoc_sdram_bankmachine7_level <= (videosoc_sdram_bankmachine7_level - 1'd1);
		end
	end
	if (videosoc_sdram_bankmachine7_wait) begin
		if ((~videosoc_sdram_bankmachine7_done)) begin
			videosoc_sdram_bankmachine7_count <= (videosoc_sdram_bankmachine7_count - 1'd1);
		end
	end else begin
		videosoc_sdram_bankmachine7_count <= 3'd5;
	end
	bankmachine7_state <= bankmachine7_next_state;
	if ((~videosoc_sdram_en0)) begin
		videosoc_sdram_time0 <= 5'd31;
	end else begin
		if ((~videosoc_sdram_max_time0)) begin
			videosoc_sdram_time0 <= (videosoc_sdram_time0 - 1'd1);
		end
	end
	if ((~videosoc_sdram_en1)) begin
		videosoc_sdram_time1 <= 4'd15;
	end else begin
		if ((~videosoc_sdram_max_time1)) begin
			videosoc_sdram_time1 <= (videosoc_sdram_time1 - 1'd1);
		end
	end
	if (videosoc_sdram_choose_cmd_ce) begin
		case (videosoc_sdram_choose_cmd_grant)
			1'd0: begin
				if (videosoc_sdram_choose_cmd_request[1]) begin
					videosoc_sdram_choose_cmd_grant <= 1'd1;
				end else begin
					if (videosoc_sdram_choose_cmd_request[2]) begin
						videosoc_sdram_choose_cmd_grant <= 2'd2;
					end else begin
						if (videosoc_sdram_choose_cmd_request[3]) begin
							videosoc_sdram_choose_cmd_grant <= 2'd3;
						end else begin
							if (videosoc_sdram_choose_cmd_request[4]) begin
								videosoc_sdram_choose_cmd_grant <= 3'd4;
							end else begin
								if (videosoc_sdram_choose_cmd_request[5]) begin
									videosoc_sdram_choose_cmd_grant <= 3'd5;
								end else begin
									if (videosoc_sdram_choose_cmd_request[6]) begin
										videosoc_sdram_choose_cmd_grant <= 3'd6;
									end else begin
										if (videosoc_sdram_choose_cmd_request[7]) begin
											videosoc_sdram_choose_cmd_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (videosoc_sdram_choose_cmd_request[2]) begin
					videosoc_sdram_choose_cmd_grant <= 2'd2;
				end else begin
					if (videosoc_sdram_choose_cmd_request[3]) begin
						videosoc_sdram_choose_cmd_grant <= 2'd3;
					end else begin
						if (videosoc_sdram_choose_cmd_request[4]) begin
							videosoc_sdram_choose_cmd_grant <= 3'd4;
						end else begin
							if (videosoc_sdram_choose_cmd_request[5]) begin
								videosoc_sdram_choose_cmd_grant <= 3'd5;
							end else begin
								if (videosoc_sdram_choose_cmd_request[6]) begin
									videosoc_sdram_choose_cmd_grant <= 3'd6;
								end else begin
									if (videosoc_sdram_choose_cmd_request[7]) begin
										videosoc_sdram_choose_cmd_grant <= 3'd7;
									end else begin
										if (videosoc_sdram_choose_cmd_request[0]) begin
											videosoc_sdram_choose_cmd_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (videosoc_sdram_choose_cmd_request[3]) begin
					videosoc_sdram_choose_cmd_grant <= 2'd3;
				end else begin
					if (videosoc_sdram_choose_cmd_request[4]) begin
						videosoc_sdram_choose_cmd_grant <= 3'd4;
					end else begin
						if (videosoc_sdram_choose_cmd_request[5]) begin
							videosoc_sdram_choose_cmd_grant <= 3'd5;
						end else begin
							if (videosoc_sdram_choose_cmd_request[6]) begin
								videosoc_sdram_choose_cmd_grant <= 3'd6;
							end else begin
								if (videosoc_sdram_choose_cmd_request[7]) begin
									videosoc_sdram_choose_cmd_grant <= 3'd7;
								end else begin
									if (videosoc_sdram_choose_cmd_request[0]) begin
										videosoc_sdram_choose_cmd_grant <= 1'd0;
									end else begin
										if (videosoc_sdram_choose_cmd_request[1]) begin
											videosoc_sdram_choose_cmd_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (videosoc_sdram_choose_cmd_request[4]) begin
					videosoc_sdram_choose_cmd_grant <= 3'd4;
				end else begin
					if (videosoc_sdram_choose_cmd_request[5]) begin
						videosoc_sdram_choose_cmd_grant <= 3'd5;
					end else begin
						if (videosoc_sdram_choose_cmd_request[6]) begin
							videosoc_sdram_choose_cmd_grant <= 3'd6;
						end else begin
							if (videosoc_sdram_choose_cmd_request[7]) begin
								videosoc_sdram_choose_cmd_grant <= 3'd7;
							end else begin
								if (videosoc_sdram_choose_cmd_request[0]) begin
									videosoc_sdram_choose_cmd_grant <= 1'd0;
								end else begin
									if (videosoc_sdram_choose_cmd_request[1]) begin
										videosoc_sdram_choose_cmd_grant <= 1'd1;
									end else begin
										if (videosoc_sdram_choose_cmd_request[2]) begin
											videosoc_sdram_choose_cmd_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (videosoc_sdram_choose_cmd_request[5]) begin
					videosoc_sdram_choose_cmd_grant <= 3'd5;
				end else begin
					if (videosoc_sdram_choose_cmd_request[6]) begin
						videosoc_sdram_choose_cmd_grant <= 3'd6;
					end else begin
						if (videosoc_sdram_choose_cmd_request[7]) begin
							videosoc_sdram_choose_cmd_grant <= 3'd7;
						end else begin
							if (videosoc_sdram_choose_cmd_request[0]) begin
								videosoc_sdram_choose_cmd_grant <= 1'd0;
							end else begin
								if (videosoc_sdram_choose_cmd_request[1]) begin
									videosoc_sdram_choose_cmd_grant <= 1'd1;
								end else begin
									if (videosoc_sdram_choose_cmd_request[2]) begin
										videosoc_sdram_choose_cmd_grant <= 2'd2;
									end else begin
										if (videosoc_sdram_choose_cmd_request[3]) begin
											videosoc_sdram_choose_cmd_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (videosoc_sdram_choose_cmd_request[6]) begin
					videosoc_sdram_choose_cmd_grant <= 3'd6;
				end else begin
					if (videosoc_sdram_choose_cmd_request[7]) begin
						videosoc_sdram_choose_cmd_grant <= 3'd7;
					end else begin
						if (videosoc_sdram_choose_cmd_request[0]) begin
							videosoc_sdram_choose_cmd_grant <= 1'd0;
						end else begin
							if (videosoc_sdram_choose_cmd_request[1]) begin
								videosoc_sdram_choose_cmd_grant <= 1'd1;
							end else begin
								if (videosoc_sdram_choose_cmd_request[2]) begin
									videosoc_sdram_choose_cmd_grant <= 2'd2;
								end else begin
									if (videosoc_sdram_choose_cmd_request[3]) begin
										videosoc_sdram_choose_cmd_grant <= 2'd3;
									end else begin
										if (videosoc_sdram_choose_cmd_request[4]) begin
											videosoc_sdram_choose_cmd_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (videosoc_sdram_choose_cmd_request[7]) begin
					videosoc_sdram_choose_cmd_grant <= 3'd7;
				end else begin
					if (videosoc_sdram_choose_cmd_request[0]) begin
						videosoc_sdram_choose_cmd_grant <= 1'd0;
					end else begin
						if (videosoc_sdram_choose_cmd_request[1]) begin
							videosoc_sdram_choose_cmd_grant <= 1'd1;
						end else begin
							if (videosoc_sdram_choose_cmd_request[2]) begin
								videosoc_sdram_choose_cmd_grant <= 2'd2;
							end else begin
								if (videosoc_sdram_choose_cmd_request[3]) begin
									videosoc_sdram_choose_cmd_grant <= 2'd3;
								end else begin
									if (videosoc_sdram_choose_cmd_request[4]) begin
										videosoc_sdram_choose_cmd_grant <= 3'd4;
									end else begin
										if (videosoc_sdram_choose_cmd_request[5]) begin
											videosoc_sdram_choose_cmd_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (videosoc_sdram_choose_cmd_request[0]) begin
					videosoc_sdram_choose_cmd_grant <= 1'd0;
				end else begin
					if (videosoc_sdram_choose_cmd_request[1]) begin
						videosoc_sdram_choose_cmd_grant <= 1'd1;
					end else begin
						if (videosoc_sdram_choose_cmd_request[2]) begin
							videosoc_sdram_choose_cmd_grant <= 2'd2;
						end else begin
							if (videosoc_sdram_choose_cmd_request[3]) begin
								videosoc_sdram_choose_cmd_grant <= 2'd3;
							end else begin
								if (videosoc_sdram_choose_cmd_request[4]) begin
									videosoc_sdram_choose_cmd_grant <= 3'd4;
								end else begin
									if (videosoc_sdram_choose_cmd_request[5]) begin
										videosoc_sdram_choose_cmd_grant <= 3'd5;
									end else begin
										if (videosoc_sdram_choose_cmd_request[6]) begin
											videosoc_sdram_choose_cmd_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (videosoc_sdram_choose_req_ce) begin
		case (videosoc_sdram_choose_req_grant)
			1'd0: begin
				if (videosoc_sdram_choose_req_request[1]) begin
					videosoc_sdram_choose_req_grant <= 1'd1;
				end else begin
					if (videosoc_sdram_choose_req_request[2]) begin
						videosoc_sdram_choose_req_grant <= 2'd2;
					end else begin
						if (videosoc_sdram_choose_req_request[3]) begin
							videosoc_sdram_choose_req_grant <= 2'd3;
						end else begin
							if (videosoc_sdram_choose_req_request[4]) begin
								videosoc_sdram_choose_req_grant <= 3'd4;
							end else begin
								if (videosoc_sdram_choose_req_request[5]) begin
									videosoc_sdram_choose_req_grant <= 3'd5;
								end else begin
									if (videosoc_sdram_choose_req_request[6]) begin
										videosoc_sdram_choose_req_grant <= 3'd6;
									end else begin
										if (videosoc_sdram_choose_req_request[7]) begin
											videosoc_sdram_choose_req_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (videosoc_sdram_choose_req_request[2]) begin
					videosoc_sdram_choose_req_grant <= 2'd2;
				end else begin
					if (videosoc_sdram_choose_req_request[3]) begin
						videosoc_sdram_choose_req_grant <= 2'd3;
					end else begin
						if (videosoc_sdram_choose_req_request[4]) begin
							videosoc_sdram_choose_req_grant <= 3'd4;
						end else begin
							if (videosoc_sdram_choose_req_request[5]) begin
								videosoc_sdram_choose_req_grant <= 3'd5;
							end else begin
								if (videosoc_sdram_choose_req_request[6]) begin
									videosoc_sdram_choose_req_grant <= 3'd6;
								end else begin
									if (videosoc_sdram_choose_req_request[7]) begin
										videosoc_sdram_choose_req_grant <= 3'd7;
									end else begin
										if (videosoc_sdram_choose_req_request[0]) begin
											videosoc_sdram_choose_req_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (videosoc_sdram_choose_req_request[3]) begin
					videosoc_sdram_choose_req_grant <= 2'd3;
				end else begin
					if (videosoc_sdram_choose_req_request[4]) begin
						videosoc_sdram_choose_req_grant <= 3'd4;
					end else begin
						if (videosoc_sdram_choose_req_request[5]) begin
							videosoc_sdram_choose_req_grant <= 3'd5;
						end else begin
							if (videosoc_sdram_choose_req_request[6]) begin
								videosoc_sdram_choose_req_grant <= 3'd6;
							end else begin
								if (videosoc_sdram_choose_req_request[7]) begin
									videosoc_sdram_choose_req_grant <= 3'd7;
								end else begin
									if (videosoc_sdram_choose_req_request[0]) begin
										videosoc_sdram_choose_req_grant <= 1'd0;
									end else begin
										if (videosoc_sdram_choose_req_request[1]) begin
											videosoc_sdram_choose_req_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (videosoc_sdram_choose_req_request[4]) begin
					videosoc_sdram_choose_req_grant <= 3'd4;
				end else begin
					if (videosoc_sdram_choose_req_request[5]) begin
						videosoc_sdram_choose_req_grant <= 3'd5;
					end else begin
						if (videosoc_sdram_choose_req_request[6]) begin
							videosoc_sdram_choose_req_grant <= 3'd6;
						end else begin
							if (videosoc_sdram_choose_req_request[7]) begin
								videosoc_sdram_choose_req_grant <= 3'd7;
							end else begin
								if (videosoc_sdram_choose_req_request[0]) begin
									videosoc_sdram_choose_req_grant <= 1'd0;
								end else begin
									if (videosoc_sdram_choose_req_request[1]) begin
										videosoc_sdram_choose_req_grant <= 1'd1;
									end else begin
										if (videosoc_sdram_choose_req_request[2]) begin
											videosoc_sdram_choose_req_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (videosoc_sdram_choose_req_request[5]) begin
					videosoc_sdram_choose_req_grant <= 3'd5;
				end else begin
					if (videosoc_sdram_choose_req_request[6]) begin
						videosoc_sdram_choose_req_grant <= 3'd6;
					end else begin
						if (videosoc_sdram_choose_req_request[7]) begin
							videosoc_sdram_choose_req_grant <= 3'd7;
						end else begin
							if (videosoc_sdram_choose_req_request[0]) begin
								videosoc_sdram_choose_req_grant <= 1'd0;
							end else begin
								if (videosoc_sdram_choose_req_request[1]) begin
									videosoc_sdram_choose_req_grant <= 1'd1;
								end else begin
									if (videosoc_sdram_choose_req_request[2]) begin
										videosoc_sdram_choose_req_grant <= 2'd2;
									end else begin
										if (videosoc_sdram_choose_req_request[3]) begin
											videosoc_sdram_choose_req_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (videosoc_sdram_choose_req_request[6]) begin
					videosoc_sdram_choose_req_grant <= 3'd6;
				end else begin
					if (videosoc_sdram_choose_req_request[7]) begin
						videosoc_sdram_choose_req_grant <= 3'd7;
					end else begin
						if (videosoc_sdram_choose_req_request[0]) begin
							videosoc_sdram_choose_req_grant <= 1'd0;
						end else begin
							if (videosoc_sdram_choose_req_request[1]) begin
								videosoc_sdram_choose_req_grant <= 1'd1;
							end else begin
								if (videosoc_sdram_choose_req_request[2]) begin
									videosoc_sdram_choose_req_grant <= 2'd2;
								end else begin
									if (videosoc_sdram_choose_req_request[3]) begin
										videosoc_sdram_choose_req_grant <= 2'd3;
									end else begin
										if (videosoc_sdram_choose_req_request[4]) begin
											videosoc_sdram_choose_req_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (videosoc_sdram_choose_req_request[7]) begin
					videosoc_sdram_choose_req_grant <= 3'd7;
				end else begin
					if (videosoc_sdram_choose_req_request[0]) begin
						videosoc_sdram_choose_req_grant <= 1'd0;
					end else begin
						if (videosoc_sdram_choose_req_request[1]) begin
							videosoc_sdram_choose_req_grant <= 1'd1;
						end else begin
							if (videosoc_sdram_choose_req_request[2]) begin
								videosoc_sdram_choose_req_grant <= 2'd2;
							end else begin
								if (videosoc_sdram_choose_req_request[3]) begin
									videosoc_sdram_choose_req_grant <= 2'd3;
								end else begin
									if (videosoc_sdram_choose_req_request[4]) begin
										videosoc_sdram_choose_req_grant <= 3'd4;
									end else begin
										if (videosoc_sdram_choose_req_request[5]) begin
											videosoc_sdram_choose_req_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (videosoc_sdram_choose_req_request[0]) begin
					videosoc_sdram_choose_req_grant <= 1'd0;
				end else begin
					if (videosoc_sdram_choose_req_request[1]) begin
						videosoc_sdram_choose_req_grant <= 1'd1;
					end else begin
						if (videosoc_sdram_choose_req_request[2]) begin
							videosoc_sdram_choose_req_grant <= 2'd2;
						end else begin
							if (videosoc_sdram_choose_req_request[3]) begin
								videosoc_sdram_choose_req_grant <= 2'd3;
							end else begin
								if (videosoc_sdram_choose_req_request[4]) begin
									videosoc_sdram_choose_req_grant <= 3'd4;
								end else begin
									if (videosoc_sdram_choose_req_request[5]) begin
										videosoc_sdram_choose_req_grant <= 3'd5;
									end else begin
										if (videosoc_sdram_choose_req_request[6]) begin
											videosoc_sdram_choose_req_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	videosoc_sdram_dfi_p0_address <= sync_rhs_array_muxed0;
	videosoc_sdram_dfi_p0_bank <= sync_rhs_array_muxed1;
	videosoc_sdram_dfi_p0_cas_n <= (~sync_rhs_array_muxed2);
	videosoc_sdram_dfi_p0_ras_n <= (~sync_rhs_array_muxed3);
	videosoc_sdram_dfi_p0_we_n <= (~sync_rhs_array_muxed4);
	videosoc_sdram_dfi_p0_rddata_en <= sync_rhs_array_muxed5;
	videosoc_sdram_dfi_p0_wrdata_en <= sync_rhs_array_muxed6;
	videosoc_sdram_dfi_p1_address <= sync_rhs_array_muxed7;
	videosoc_sdram_dfi_p1_bank <= sync_rhs_array_muxed8;
	videosoc_sdram_dfi_p1_cas_n <= (~sync_rhs_array_muxed9);
	videosoc_sdram_dfi_p1_ras_n <= (~sync_rhs_array_muxed10);
	videosoc_sdram_dfi_p1_we_n <= (~sync_rhs_array_muxed11);
	videosoc_sdram_dfi_p1_rddata_en <= sync_rhs_array_muxed12;
	videosoc_sdram_dfi_p1_wrdata_en <= sync_rhs_array_muxed13;
	videosoc_sdram_dfi_p2_address <= sync_rhs_array_muxed14;
	videosoc_sdram_dfi_p2_bank <= sync_rhs_array_muxed15;
	videosoc_sdram_dfi_p2_cas_n <= (~sync_rhs_array_muxed16);
	videosoc_sdram_dfi_p2_ras_n <= (~sync_rhs_array_muxed17);
	videosoc_sdram_dfi_p2_we_n <= (~sync_rhs_array_muxed18);
	videosoc_sdram_dfi_p2_rddata_en <= sync_rhs_array_muxed19;
	videosoc_sdram_dfi_p2_wrdata_en <= sync_rhs_array_muxed20;
	videosoc_sdram_dfi_p3_address <= sync_rhs_array_muxed21;
	videosoc_sdram_dfi_p3_bank <= sync_rhs_array_muxed22;
	videosoc_sdram_dfi_p3_cas_n <= (~sync_rhs_array_muxed23);
	videosoc_sdram_dfi_p3_ras_n <= (~sync_rhs_array_muxed24);
	videosoc_sdram_dfi_p3_we_n <= (~sync_rhs_array_muxed25);
	videosoc_sdram_dfi_p3_rddata_en <= sync_rhs_array_muxed26;
	videosoc_sdram_dfi_p3_wrdata_en <= sync_rhs_array_muxed27;
	multiplexer_state <= multiplexer_next_state;
	videosoc_sdram_bandwidth_cmd_valid <= videosoc_sdram_choose_req_cmd_valid;
	videosoc_sdram_bandwidth_cmd_ready <= videosoc_sdram_choose_req_cmd_ready;
	videosoc_sdram_bandwidth_cmd_is_read <= videosoc_sdram_choose_req_cmd_payload_is_read;
	videosoc_sdram_bandwidth_cmd_is_write <= videosoc_sdram_choose_req_cmd_payload_is_write;
	{videosoc_sdram_bandwidth_period, videosoc_sdram_bandwidth_counter} <= (videosoc_sdram_bandwidth_counter + 1'd1);
	if (videosoc_sdram_bandwidth_period) begin
		videosoc_sdram_bandwidth_nreads_r <= videosoc_sdram_bandwidth_nreads;
		videosoc_sdram_bandwidth_nwrites_r <= videosoc_sdram_bandwidth_nwrites;
		videosoc_sdram_bandwidth_nreads <= 1'd0;
		videosoc_sdram_bandwidth_nwrites <= 1'd0;
	end else begin
		if ((videosoc_sdram_bandwidth_cmd_valid & videosoc_sdram_bandwidth_cmd_ready)) begin
			if (videosoc_sdram_bandwidth_cmd_is_read) begin
				videosoc_sdram_bandwidth_nreads <= (videosoc_sdram_bandwidth_nreads + 1'd1);
			end
			if (videosoc_sdram_bandwidth_cmd_is_write) begin
				videosoc_sdram_bandwidth_nwrites <= (videosoc_sdram_bandwidth_nwrites + 1'd1);
			end
		end
	end
	if (videosoc_sdram_bandwidth_update_re) begin
		videosoc_sdram_bandwidth_nreads_status <= videosoc_sdram_bandwidth_nreads_r;
		videosoc_sdram_bandwidth_nwrites_status <= videosoc_sdram_bandwidth_nwrites_r;
	end
	new_master_wdata_ready0 <= ((((((((1'd0 | ((roundrobin0_grant == 1'd0) & videosoc_sdram_interface_bank0_wdata_ready)) | ((roundrobin1_grant == 1'd0) & videosoc_sdram_interface_bank1_wdata_ready)) | ((roundrobin2_grant == 1'd0) & videosoc_sdram_interface_bank2_wdata_ready)) | ((roundrobin3_grant == 1'd0) & videosoc_sdram_interface_bank3_wdata_ready)) | ((roundrobin4_grant == 1'd0) & videosoc_sdram_interface_bank4_wdata_ready)) | ((roundrobin5_grant == 1'd0) & videosoc_sdram_interface_bank5_wdata_ready)) | ((roundrobin6_grant == 1'd0) & videosoc_sdram_interface_bank6_wdata_ready)) | ((roundrobin7_grant == 1'd0) & videosoc_sdram_interface_bank7_wdata_ready));
	new_master_wdata_ready1 <= new_master_wdata_ready0;
	new_master_wdata_ready2 <= new_master_wdata_ready1;
	new_master_wdata_ready3 <= ((((((((1'd0 | ((roundrobin0_grant == 1'd1) & videosoc_sdram_interface_bank0_wdata_ready)) | ((roundrobin1_grant == 1'd1) & videosoc_sdram_interface_bank1_wdata_ready)) | ((roundrobin2_grant == 1'd1) & videosoc_sdram_interface_bank2_wdata_ready)) | ((roundrobin3_grant == 1'd1) & videosoc_sdram_interface_bank3_wdata_ready)) | ((roundrobin4_grant == 1'd1) & videosoc_sdram_interface_bank4_wdata_ready)) | ((roundrobin5_grant == 1'd1) & videosoc_sdram_interface_bank5_wdata_ready)) | ((roundrobin6_grant == 1'd1) & videosoc_sdram_interface_bank6_wdata_ready)) | ((roundrobin7_grant == 1'd1) & videosoc_sdram_interface_bank7_wdata_ready));
	new_master_wdata_ready4 <= new_master_wdata_ready3;
	new_master_wdata_ready5 <= new_master_wdata_ready4;
	new_master_wdata_ready6 <= ((((((((1'd0 | ((roundrobin0_grant == 2'd2) & videosoc_sdram_interface_bank0_wdata_ready)) | ((roundrobin1_grant == 2'd2) & videosoc_sdram_interface_bank1_wdata_ready)) | ((roundrobin2_grant == 2'd2) & videosoc_sdram_interface_bank2_wdata_ready)) | ((roundrobin3_grant == 2'd2) & videosoc_sdram_interface_bank3_wdata_ready)) | ((roundrobin4_grant == 2'd2) & videosoc_sdram_interface_bank4_wdata_ready)) | ((roundrobin5_grant == 2'd2) & videosoc_sdram_interface_bank5_wdata_ready)) | ((roundrobin6_grant == 2'd2) & videosoc_sdram_interface_bank6_wdata_ready)) | ((roundrobin7_grant == 2'd2) & videosoc_sdram_interface_bank7_wdata_ready));
	new_master_wdata_ready7 <= new_master_wdata_ready6;
	new_master_wdata_ready8 <= new_master_wdata_ready7;
	new_master_rdata_valid0 <= ((((((((1'd0 | ((roundrobin0_grant == 1'd0) & videosoc_sdram_interface_bank0_rdata_valid)) | ((roundrobin1_grant == 1'd0) & videosoc_sdram_interface_bank1_rdata_valid)) | ((roundrobin2_grant == 1'd0) & videosoc_sdram_interface_bank2_rdata_valid)) | ((roundrobin3_grant == 1'd0) & videosoc_sdram_interface_bank3_rdata_valid)) | ((roundrobin4_grant == 1'd0) & videosoc_sdram_interface_bank4_rdata_valid)) | ((roundrobin5_grant == 1'd0) & videosoc_sdram_interface_bank5_rdata_valid)) | ((roundrobin6_grant == 1'd0) & videosoc_sdram_interface_bank6_rdata_valid)) | ((roundrobin7_grant == 1'd0) & videosoc_sdram_interface_bank7_rdata_valid));
	new_master_rdata_valid1 <= new_master_rdata_valid0;
	new_master_rdata_valid2 <= new_master_rdata_valid1;
	new_master_rdata_valid3 <= new_master_rdata_valid2;
	new_master_rdata_valid4 <= new_master_rdata_valid3;
	new_master_rdata_valid5 <= new_master_rdata_valid4;
	new_master_rdata_valid6 <= new_master_rdata_valid5;
	new_master_rdata_valid7 <= ((((((((1'd0 | ((roundrobin0_grant == 1'd1) & videosoc_sdram_interface_bank0_rdata_valid)) | ((roundrobin1_grant == 1'd1) & videosoc_sdram_interface_bank1_rdata_valid)) | ((roundrobin2_grant == 1'd1) & videosoc_sdram_interface_bank2_rdata_valid)) | ((roundrobin3_grant == 1'd1) & videosoc_sdram_interface_bank3_rdata_valid)) | ((roundrobin4_grant == 1'd1) & videosoc_sdram_interface_bank4_rdata_valid)) | ((roundrobin5_grant == 1'd1) & videosoc_sdram_interface_bank5_rdata_valid)) | ((roundrobin6_grant == 1'd1) & videosoc_sdram_interface_bank6_rdata_valid)) | ((roundrobin7_grant == 1'd1) & videosoc_sdram_interface_bank7_rdata_valid));
	new_master_rdata_valid8 <= new_master_rdata_valid7;
	new_master_rdata_valid9 <= new_master_rdata_valid8;
	new_master_rdata_valid10 <= new_master_rdata_valid9;
	new_master_rdata_valid11 <= new_master_rdata_valid10;
	new_master_rdata_valid12 <= new_master_rdata_valid11;
	new_master_rdata_valid13 <= new_master_rdata_valid12;
	new_master_rdata_valid14 <= ((((((((1'd0 | ((roundrobin0_grant == 2'd2) & videosoc_sdram_interface_bank0_rdata_valid)) | ((roundrobin1_grant == 2'd2) & videosoc_sdram_interface_bank1_rdata_valid)) | ((roundrobin2_grant == 2'd2) & videosoc_sdram_interface_bank2_rdata_valid)) | ((roundrobin3_grant == 2'd2) & videosoc_sdram_interface_bank3_rdata_valid)) | ((roundrobin4_grant == 2'd2) & videosoc_sdram_interface_bank4_rdata_valid)) | ((roundrobin5_grant == 2'd2) & videosoc_sdram_interface_bank5_rdata_valid)) | ((roundrobin6_grant == 2'd2) & videosoc_sdram_interface_bank6_rdata_valid)) | ((roundrobin7_grant == 2'd2) & videosoc_sdram_interface_bank7_rdata_valid));
	new_master_rdata_valid15 <= new_master_rdata_valid14;
	new_master_rdata_valid16 <= new_master_rdata_valid15;
	new_master_rdata_valid17 <= new_master_rdata_valid16;
	new_master_rdata_valid18 <= new_master_rdata_valid17;
	new_master_rdata_valid19 <= new_master_rdata_valid18;
	new_master_rdata_valid20 <= new_master_rdata_valid19;
	hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary <= hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary;
	hdmi_out0_dram_port_cmd_fifo_graycounter1_q <= hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next;
	hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary <= hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary;
	hdmi_out0_dram_port_rdata_fifo_graycounter0_q <= hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next;
	if (roundrobin0_ce) begin
		case (roundrobin0_grant)
			1'd0: begin
				if (roundrobin0_request[1]) begin
					roundrobin0_grant <= 1'd1;
				end else begin
					if (roundrobin0_request[2]) begin
						roundrobin0_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin0_request[2]) begin
					roundrobin0_grant <= 2'd2;
				end else begin
					if (roundrobin0_request[0]) begin
						roundrobin0_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin0_request[0]) begin
					roundrobin0_grant <= 1'd0;
				end else begin
					if (roundrobin0_request[1]) begin
						roundrobin0_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (roundrobin1_ce) begin
		case (roundrobin1_grant)
			1'd0: begin
				if (roundrobin1_request[1]) begin
					roundrobin1_grant <= 1'd1;
				end else begin
					if (roundrobin1_request[2]) begin
						roundrobin1_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin1_request[2]) begin
					roundrobin1_grant <= 2'd2;
				end else begin
					if (roundrobin1_request[0]) begin
						roundrobin1_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin1_request[0]) begin
					roundrobin1_grant <= 1'd0;
				end else begin
					if (roundrobin1_request[1]) begin
						roundrobin1_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (roundrobin2_ce) begin
		case (roundrobin2_grant)
			1'd0: begin
				if (roundrobin2_request[1]) begin
					roundrobin2_grant <= 1'd1;
				end else begin
					if (roundrobin2_request[2]) begin
						roundrobin2_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin2_request[2]) begin
					roundrobin2_grant <= 2'd2;
				end else begin
					if (roundrobin2_request[0]) begin
						roundrobin2_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin2_request[0]) begin
					roundrobin2_grant <= 1'd0;
				end else begin
					if (roundrobin2_request[1]) begin
						roundrobin2_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (roundrobin3_ce) begin
		case (roundrobin3_grant)
			1'd0: begin
				if (roundrobin3_request[1]) begin
					roundrobin3_grant <= 1'd1;
				end else begin
					if (roundrobin3_request[2]) begin
						roundrobin3_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin3_request[2]) begin
					roundrobin3_grant <= 2'd2;
				end else begin
					if (roundrobin3_request[0]) begin
						roundrobin3_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin3_request[0]) begin
					roundrobin3_grant <= 1'd0;
				end else begin
					if (roundrobin3_request[1]) begin
						roundrobin3_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (roundrobin4_ce) begin
		case (roundrobin4_grant)
			1'd0: begin
				if (roundrobin4_request[1]) begin
					roundrobin4_grant <= 1'd1;
				end else begin
					if (roundrobin4_request[2]) begin
						roundrobin4_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin4_request[2]) begin
					roundrobin4_grant <= 2'd2;
				end else begin
					if (roundrobin4_request[0]) begin
						roundrobin4_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin4_request[0]) begin
					roundrobin4_grant <= 1'd0;
				end else begin
					if (roundrobin4_request[1]) begin
						roundrobin4_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (roundrobin5_ce) begin
		case (roundrobin5_grant)
			1'd0: begin
				if (roundrobin5_request[1]) begin
					roundrobin5_grant <= 1'd1;
				end else begin
					if (roundrobin5_request[2]) begin
						roundrobin5_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin5_request[2]) begin
					roundrobin5_grant <= 2'd2;
				end else begin
					if (roundrobin5_request[0]) begin
						roundrobin5_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin5_request[0]) begin
					roundrobin5_grant <= 1'd0;
				end else begin
					if (roundrobin5_request[1]) begin
						roundrobin5_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (roundrobin6_ce) begin
		case (roundrobin6_grant)
			1'd0: begin
				if (roundrobin6_request[1]) begin
					roundrobin6_grant <= 1'd1;
				end else begin
					if (roundrobin6_request[2]) begin
						roundrobin6_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin6_request[2]) begin
					roundrobin6_grant <= 2'd2;
				end else begin
					if (roundrobin6_request[0]) begin
						roundrobin6_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin6_request[0]) begin
					roundrobin6_grant <= 1'd0;
				end else begin
					if (roundrobin6_request[1]) begin
						roundrobin6_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (roundrobin7_ce) begin
		case (roundrobin7_grant)
			1'd0: begin
				if (roundrobin7_request[1]) begin
					roundrobin7_grant <= 1'd1;
				end else begin
					if (roundrobin7_request[2]) begin
						roundrobin7_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (roundrobin7_request[2]) begin
					roundrobin7_grant <= 2'd2;
				end else begin
					if (roundrobin7_request[0]) begin
						roundrobin7_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (roundrobin7_request[0]) begin
					roundrobin7_grant <= 1'd0;
				end else begin
					if (roundrobin7_request[1]) begin
						roundrobin7_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	videosoc_adr_offset_r <= videosoc_interface0_wb_sdram_adr[1:0];
	fullmemorywe_state <= fullmemorywe_next_state;
	litedramwishbonebridge_state <= litedramwishbonebridge_next_state;
	if ((videosoc_i == 1'd0)) begin
		videosoc_clk1 <= 1'd1;
		videosoc_miso <= spiflash_1x_miso;
	end
	if ((videosoc_i == 1'd1)) begin
		videosoc_i <= 1'd0;
		videosoc_clk1 <= 1'd0;
		videosoc_sr <= {videosoc_sr[30:0], videosoc_miso};
	end else begin
		videosoc_i <= (videosoc_i + 1'd1);
	end
	if ((((videosoc_bus_cyc & videosoc_bus_stb) & (videosoc_i == 1'd1)) & (videosoc_counter == 1'd0))) begin
		videosoc_cs_n <= 1'd0;
		videosoc_sr[31:24] <= 4'd11;
	end
	if ((videosoc_counter == 5'd16)) begin
		videosoc_sr[31:8] <= {videosoc_bus_adr, {2{1'd0}}};
	end
	if ((videosoc_counter == 7'd64)) begin
	end
	if ((videosoc_counter == 8'd146)) begin
		videosoc_bus_ack <= 1'd1;
		videosoc_cs_n <= 1'd1;
	end
	if ((videosoc_counter == 8'd147)) begin
		videosoc_bus_ack <= 1'd0;
	end
	if ((videosoc_counter == 8'd149)) begin
	end
	if ((videosoc_counter == 8'd149)) begin
		videosoc_counter <= 1'd0;
	end else begin
		if ((videosoc_counter != 1'd0)) begin
			videosoc_counter <= (videosoc_counter + 1'd1);
		end else begin
			if (((videosoc_bus_cyc & videosoc_bus_stb) & (videosoc_i == 1'd1))) begin
				videosoc_counter <= 1'd1;
			end
		end
	end
	if (ethphy_counter_ce) begin
		ethphy_counter <= (ethphy_counter + 1'd1);
	end
	if (ethmac_ps_preamble_error_o) begin
		ethmac_preamble_errors_status <= (ethmac_preamble_errors_status + 1'd1);
	end
	if (ethmac_ps_crc_error_o) begin
		ethmac_crc_errors_status <= (ethmac_crc_errors_status + 1'd1);
	end
	ethmac_ps_preamble_error_toggle_o_r <= ethmac_ps_preamble_error_toggle_o;
	ethmac_ps_crc_error_toggle_o_r <= ethmac_ps_crc_error_toggle_o;
	ethmac_tx_cdc_graycounter0_q_binary <= ethmac_tx_cdc_graycounter0_q_next_binary;
	ethmac_tx_cdc_graycounter0_q <= ethmac_tx_cdc_graycounter0_q_next;
	ethmac_rx_cdc_graycounter1_q_binary <= ethmac_rx_cdc_graycounter1_q_next_binary;
	ethmac_rx_cdc_graycounter1_q <= ethmac_rx_cdc_graycounter1_q_next;
	if (ethmac_writer_counter_reset) begin
		ethmac_writer_counter <= 1'd0;
	end else begin
		if (ethmac_writer_counter_ce) begin
			ethmac_writer_counter <= (ethmac_writer_counter + ethmac_writer_increment);
		end
	end
	if (ethmac_writer_slot_ce) begin
		ethmac_writer_slot <= (ethmac_writer_slot + 1'd1);
	end
	if (((ethmac_writer_fifo_syncfifo_we & ethmac_writer_fifo_syncfifo_writable) & (~ethmac_writer_fifo_replace))) begin
		ethmac_writer_fifo_produce <= (ethmac_writer_fifo_produce + 1'd1);
	end
	if (ethmac_writer_fifo_do_read) begin
		ethmac_writer_fifo_consume <= (ethmac_writer_fifo_consume + 1'd1);
	end
	if (((ethmac_writer_fifo_syncfifo_we & ethmac_writer_fifo_syncfifo_writable) & (~ethmac_writer_fifo_replace))) begin
		if ((~ethmac_writer_fifo_do_read)) begin
			ethmac_writer_fifo_level <= (ethmac_writer_fifo_level + 1'd1);
		end
	end else begin
		if (ethmac_writer_fifo_do_read) begin
			ethmac_writer_fifo_level <= (ethmac_writer_fifo_level - 1'd1);
		end
	end
	liteethmacsramwriter_state <= liteethmacsramwriter_next_state;
	if (ethmac_writer_errors_status_liteethmac_next_value_ce) begin
		ethmac_writer_errors_status <= ethmac_writer_errors_status_liteethmac_next_value;
	end
	if (ethmac_reader_counter_reset) begin
		ethmac_reader_counter <= 1'd0;
	end else begin
		if (ethmac_reader_counter_ce) begin
			ethmac_reader_counter <= (ethmac_reader_counter + 3'd4);
		end
	end
	ethmac_reader_last_d <= ethmac_reader_last;
	if (ethmac_reader_done_clear) begin
		ethmac_reader_done_pending <= 1'd0;
	end
	if (ethmac_reader_done_trigger) begin
		ethmac_reader_done_pending <= 1'd1;
	end
	if (((ethmac_reader_fifo_syncfifo_we & ethmac_reader_fifo_syncfifo_writable) & (~ethmac_reader_fifo_replace))) begin
		ethmac_reader_fifo_produce <= (ethmac_reader_fifo_produce + 1'd1);
	end
	if (ethmac_reader_fifo_do_read) begin
		ethmac_reader_fifo_consume <= (ethmac_reader_fifo_consume + 1'd1);
	end
	if (((ethmac_reader_fifo_syncfifo_we & ethmac_reader_fifo_syncfifo_writable) & (~ethmac_reader_fifo_replace))) begin
		if ((~ethmac_reader_fifo_do_read)) begin
			ethmac_reader_fifo_level <= (ethmac_reader_fifo_level + 1'd1);
		end
	end else begin
		if (ethmac_reader_fifo_do_read) begin
			ethmac_reader_fifo_level <= (ethmac_reader_fifo_level - 1'd1);
		end
	end
	liteethmacsramreader_state <= liteethmacsramreader_next_state;
	ethmac_sram0_bus_ack0 <= 1'd0;
	if (((ethmac_sram0_bus_cyc0 & ethmac_sram0_bus_stb0) & (~ethmac_sram0_bus_ack0))) begin
		ethmac_sram0_bus_ack0 <= 1'd1;
	end
	ethmac_sram1_bus_ack0 <= 1'd0;
	if (((ethmac_sram1_bus_cyc0 & ethmac_sram1_bus_stb0) & (~ethmac_sram1_bus_ack0))) begin
		ethmac_sram1_bus_ack0 <= 1'd1;
	end
	ethmac_sram0_bus_ack1 <= 1'd0;
	if (((ethmac_sram0_bus_cyc1 & ethmac_sram0_bus_stb1) & (~ethmac_sram0_bus_ack1))) begin
		ethmac_sram0_bus_ack1 <= 1'd1;
	end
	ethmac_sram1_bus_ack1 <= 1'd0;
	if (((ethmac_sram1_bus_cyc1 & ethmac_sram1_bus_stb1) & (~ethmac_sram1_bus_ack1))) begin
		ethmac_sram1_bus_ack1 <= 1'd1;
	end
	ethmac_slave_sel_r <= ethmac_slave_sel;
	edid_sda_drv_reg <= edid_sda_drv;
	{edid_samp_carry, edid_samp_count} <= (edid_samp_count + 1'd1);
	if (edid_samp_carry) begin
		edid_scl_i <= edid_scl_raw;
		edid_sda_i <= edid_sda_raw;
	end
	edid_scl_r <= edid_scl_i;
	edid_sda_r <= edid_sda_i;
	if (edid_start) begin
		edid_counter <= 1'd0;
	end
	if (edid_scl_rising) begin
		if ((edid_counter == 4'd8)) begin
			edid_counter <= 1'd0;
		end else begin
			edid_counter <= (edid_counter + 1'd1);
			edid_din <= {edid_din[6:0], edid_sda_i};
		end
	end
	if (edid_update_is_read) begin
		edid_is_read <= edid_din[0];
	end
	if (edid_oc_load) begin
		edid_offset_counter <= edid_din;
	end else begin
		if (edid_oc_inc) begin
			edid_offset_counter <= (edid_offset_counter + 1'd1);
		end
	end
	if (edid_data_drv_en) begin
		edid_data_drv <= 1'd1;
	end else begin
		if (edid_data_drv_stop) begin
			edid_data_drv <= 1'd0;
		end
	end
	if (edid_data_drv_en) begin
		case (edid_counter)
			1'd0: begin
				edid_data_bit <= edid_dat_r[7];
			end
			1'd1: begin
				edid_data_bit <= edid_dat_r[6];
			end
			2'd2: begin
				edid_data_bit <= edid_dat_r[5];
			end
			2'd3: begin
				edid_data_bit <= edid_dat_r[4];
			end
			3'd4: begin
				edid_data_bit <= edid_dat_r[3];
			end
			3'd5: begin
				edid_data_bit <= edid_dat_r[2];
			end
			3'd6: begin
				edid_data_bit <= edid_dat_r[1];
			end
			default: begin
				edid_data_bit <= edid_dat_r[0];
			end
		endcase
	end
	edid_state <= edid_next_state;
	if ((mmcm_read_re | mmcm_write_re)) begin
		mmcm_drdy_status <= 1'd0;
	end else begin
		if (mmcm_drdy) begin
			mmcm_drdy_status <= 1'd1;
		end
	end
	if (s7datacapture0_do_delay_rst_i) begin
		s7datacapture0_do_delay_rst_toggle_i <= (~s7datacapture0_do_delay_rst_toggle_i);
	end
	if (s7datacapture0_do_delay_master_inc_i) begin
		s7datacapture0_do_delay_master_inc_toggle_i <= (~s7datacapture0_do_delay_master_inc_toggle_i);
	end
	if (s7datacapture0_do_delay_master_dec_i) begin
		s7datacapture0_do_delay_master_dec_toggle_i <= (~s7datacapture0_do_delay_master_dec_toggle_i);
	end
	if (s7datacapture0_do_delay_slave_inc_i) begin
		s7datacapture0_do_delay_slave_inc_toggle_i <= (~s7datacapture0_do_delay_slave_inc_toggle_i);
	end
	if (s7datacapture0_do_delay_slave_dec_i) begin
		s7datacapture0_do_delay_slave_dec_toggle_i <= (~s7datacapture0_do_delay_slave_dec_toggle_i);
	end
	if (s7datacapture0_do_reset_lateness_i) begin
		s7datacapture0_do_reset_lateness_toggle_i <= (~s7datacapture0_do_reset_lateness_toggle_i);
	end
	if (wer0_o) begin
		wer0_wer_counter_sys <= wer0_wer_counter_r;
	end
	if (wer0_update_re) begin
		wer0_status <= wer0_wer_counter_sys;
	end
	wer0_toggle_o_r <= wer0_toggle_o;
	if (s7datacapture1_do_delay_rst_i) begin
		s7datacapture1_do_delay_rst_toggle_i <= (~s7datacapture1_do_delay_rst_toggle_i);
	end
	if (s7datacapture1_do_delay_master_inc_i) begin
		s7datacapture1_do_delay_master_inc_toggle_i <= (~s7datacapture1_do_delay_master_inc_toggle_i);
	end
	if (s7datacapture1_do_delay_master_dec_i) begin
		s7datacapture1_do_delay_master_dec_toggle_i <= (~s7datacapture1_do_delay_master_dec_toggle_i);
	end
	if (s7datacapture1_do_delay_slave_inc_i) begin
		s7datacapture1_do_delay_slave_inc_toggle_i <= (~s7datacapture1_do_delay_slave_inc_toggle_i);
	end
	if (s7datacapture1_do_delay_slave_dec_i) begin
		s7datacapture1_do_delay_slave_dec_toggle_i <= (~s7datacapture1_do_delay_slave_dec_toggle_i);
	end
	if (s7datacapture1_do_reset_lateness_i) begin
		s7datacapture1_do_reset_lateness_toggle_i <= (~s7datacapture1_do_reset_lateness_toggle_i);
	end
	if (wer1_o) begin
		wer1_wer_counter_sys <= wer1_wer_counter_r;
	end
	if (wer1_update_re) begin
		wer1_status <= wer1_wer_counter_sys;
	end
	wer1_toggle_o_r <= wer1_toggle_o;
	if (s7datacapture2_do_delay_rst_i) begin
		s7datacapture2_do_delay_rst_toggle_i <= (~s7datacapture2_do_delay_rst_toggle_i);
	end
	if (s7datacapture2_do_delay_master_inc_i) begin
		s7datacapture2_do_delay_master_inc_toggle_i <= (~s7datacapture2_do_delay_master_inc_toggle_i);
	end
	if (s7datacapture2_do_delay_master_dec_i) begin
		s7datacapture2_do_delay_master_dec_toggle_i <= (~s7datacapture2_do_delay_master_dec_toggle_i);
	end
	if (s7datacapture2_do_delay_slave_inc_i) begin
		s7datacapture2_do_delay_slave_inc_toggle_i <= (~s7datacapture2_do_delay_slave_inc_toggle_i);
	end
	if (s7datacapture2_do_delay_slave_dec_i) begin
		s7datacapture2_do_delay_slave_dec_toggle_i <= (~s7datacapture2_do_delay_slave_dec_toggle_i);
	end
	if (s7datacapture2_do_reset_lateness_i) begin
		s7datacapture2_do_reset_lateness_toggle_i <= (~s7datacapture2_do_reset_lateness_toggle_i);
	end
	if (wer2_o) begin
		wer2_wer_counter_sys <= wer2_wer_counter_r;
	end
	if (wer2_update_re) begin
		wer2_status <= wer2_wer_counter_sys;
	end
	wer2_toggle_o_r <= wer2_toggle_o;
	if (frame_overflow_re) begin
		frame_overflow_mask <= 1'd1;
	end else begin
		if (frame_overflow_reset_ack_o) begin
			frame_overflow_mask <= 1'd0;
		end
	end
	frame_fifo_graycounter1_q_binary <= frame_fifo_graycounter1_q_next_binary;
	frame_fifo_graycounter1_q <= frame_fifo_graycounter1_q_next;
	if (frame_overflow_reset_i) begin
		frame_overflow_reset_toggle_i <= (~frame_overflow_reset_toggle_i);
	end
	frame_overflow_reset_ack_toggle_o_r <= frame_overflow_reset_ack_toggle_o;
	if (dma_reset_words) begin
		dma_current_address <= dma_slot_array_address;
		dma_mwords_remaining <= dma_frame_size_storage;
	end else begin
		if (dma_count_word) begin
			dma_current_address <= (dma_current_address + 1'd1);
			dma_mwords_remaining <= (dma_mwords_remaining - 1'd1);
		end
	end
	if (dma_slot_array_change_slot) begin
		if (dma_slot_array_slot1_address_valid) begin
			dma_slot_array_current_slot <= 1'd1;
		end
		if (dma_slot_array_slot0_address_valid) begin
			dma_slot_array_current_slot <= 1'd0;
		end
	end
	if (((dma_fifo_syncfifo_we & dma_fifo_syncfifo_writable) & (~dma_fifo_replace))) begin
		dma_fifo_produce <= (dma_fifo_produce + 1'd1);
	end
	if (dma_fifo_do_read) begin
		dma_fifo_consume <= (dma_fifo_consume + 1'd1);
	end
	if (((dma_fifo_syncfifo_we & dma_fifo_syncfifo_writable) & (~dma_fifo_replace))) begin
		if ((~dma_fifo_do_read)) begin
			dma_fifo_level <= (dma_fifo_level + 1'd1);
		end
	end else begin
		if (dma_fifo_do_read) begin
			dma_fifo_level <= (dma_fifo_level - 1'd1);
		end
	end
	dma_state <= dma_next_state;
	if (hdmi_in0_freq_period_done) begin
		hdmi_in0_freq_period_counter <= 1'd0;
	end else begin
		hdmi_in0_freq_period_counter <= (hdmi_in0_freq_period_counter + 1'd1);
	end
	hdmi_in0_freq_gray_decoder_o <= hdmi_in0_freq_gray_decoder_o_comb;
	hdmi_in0_freq_sampler_i_d <= hdmi_in0_freq_sampler_i;
	if (hdmi_in0_freq_sampler_latch) begin
		hdmi_in0_freq_sampler_counter <= 1'd0;
		hdmi_in0_freq_sampler_o <= hdmi_in0_freq_sampler_counter;
	end else begin
		hdmi_in0_freq_sampler_counter <= (hdmi_in0_freq_sampler_counter + hdmi_in0_freq_sampler_inc);
	end
	hdmi_out0_core_initiator_cdc_graycounter0_q_binary <= hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary;
	hdmi_out0_core_initiator_cdc_graycounter0_q <= hdmi_out0_core_initiator_cdc_graycounter0_q_next;
	if (hdmi_out0_core_i) begin
		hdmi_out0_core_toggle_i <= (~hdmi_out0_core_toggle_i);
	end
	if ((hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re | hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re)) begin
		hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status <= 1'd0;
	end else begin
		if (hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy) begin
			hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status <= 1'd1;
		end
	end
	case (videosoc_grant)
		1'd0: begin
			if ((~videosoc_request[0])) begin
				if (videosoc_request[1]) begin
					videosoc_grant <= 1'd1;
				end else begin
					if (videosoc_request[2]) begin
						videosoc_grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~videosoc_request[1])) begin
				if (videosoc_request[2]) begin
					videosoc_grant <= 2'd2;
				end else begin
					if (videosoc_request[0]) begin
						videosoc_grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~videosoc_request[2])) begin
				if (videosoc_request[0]) begin
					videosoc_grant <= 1'd0;
				end else begin
					if (videosoc_request[1]) begin
						videosoc_grant <= 1'd1;
					end
				end
			end
		end
	endcase
	videosoc_slave_sel_r <= videosoc_slave_sel;
	videosoc_interface0_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank0_sel) begin
		case (videosoc_interface0_bank_bus_adr[1:0])
			1'd0: begin
				videosoc_interface0_bank_bus_dat_r <= videosoc_csrbank0_dly_sel0_w;
			end
			1'd1: begin
				videosoc_interface0_bank_bus_dat_r <= videosoc_ddrphy_rdly_dq_rst_w;
			end
			2'd2: begin
				videosoc_interface0_bank_bus_dat_r <= videosoc_ddrphy_rdly_dq_inc_w;
			end
			2'd3: begin
				videosoc_interface0_bank_bus_dat_r <= videosoc_ddrphy_rdly_dq_bitslip_w;
			end
		endcase
	end
	if (videosoc_csrbank0_dly_sel0_re) begin
		videosoc_ddrphy_storage_full[1:0] <= videosoc_csrbank0_dly_sel0_r;
	end
	videosoc_ddrphy_re <= videosoc_csrbank0_dly_sel0_re;
	videosoc_interface1_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank1_sel) begin
		case (videosoc_interface1_bank_bus_adr[4:0])
			1'd0: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_slot_w;
			end
			1'd1: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_length3_w;
			end
			2'd2: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_length2_w;
			end
			2'd3: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_length1_w;
			end
			3'd4: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_length0_w;
			end
			3'd5: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_errors3_w;
			end
			3'd6: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_errors2_w;
			end
			3'd7: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_errors1_w;
			end
			4'd8: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_errors0_w;
			end
			4'd9: begin
				videosoc_interface1_bank_bus_dat_r <= ethmac_writer_status_w;
			end
			4'd10: begin
				videosoc_interface1_bank_bus_dat_r <= ethmac_writer_pending_w;
			end
			4'd11: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_writer_ev_enable0_w;
			end
			4'd12: begin
				videosoc_interface1_bank_bus_dat_r <= ethmac_reader_start_w;
			end
			4'd13: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_reader_ready_w;
			end
			4'd14: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_reader_level_w;
			end
			4'd15: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_reader_slot0_w;
			end
			5'd16: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_reader_length1_w;
			end
			5'd17: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_reader_length0_w;
			end
			5'd18: begin
				videosoc_interface1_bank_bus_dat_r <= ethmac_reader_eventmanager_status_w;
			end
			5'd19: begin
				videosoc_interface1_bank_bus_dat_r <= ethmac_reader_eventmanager_pending_w;
			end
			5'd20: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_sram_reader_ev_enable0_w;
			end
			5'd21: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_preamble_crc_w;
			end
			5'd22: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_preamble_errors3_w;
			end
			5'd23: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_preamble_errors2_w;
			end
			5'd24: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_preamble_errors1_w;
			end
			5'd25: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_preamble_errors0_w;
			end
			5'd26: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_crc_errors3_w;
			end
			5'd27: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_crc_errors2_w;
			end
			5'd28: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_crc_errors1_w;
			end
			5'd29: begin
				videosoc_interface1_bank_bus_dat_r <= videosoc_csrbank1_crc_errors0_w;
			end
		endcase
	end
	if (videosoc_csrbank1_sram_writer_ev_enable0_re) begin
		ethmac_writer_storage_full <= videosoc_csrbank1_sram_writer_ev_enable0_r;
	end
	ethmac_writer_re <= videosoc_csrbank1_sram_writer_ev_enable0_re;
	if (videosoc_csrbank1_sram_reader_slot0_re) begin
		ethmac_reader_slot_storage_full <= videosoc_csrbank1_sram_reader_slot0_r;
	end
	ethmac_reader_slot_re <= videosoc_csrbank1_sram_reader_slot0_re;
	if (videosoc_csrbank1_sram_reader_length1_re) begin
		ethmac_reader_length_storage_full[10:8] <= videosoc_csrbank1_sram_reader_length1_r;
	end
	if (videosoc_csrbank1_sram_reader_length0_re) begin
		ethmac_reader_length_storage_full[7:0] <= videosoc_csrbank1_sram_reader_length0_r;
	end
	ethmac_reader_length_re <= videosoc_csrbank1_sram_reader_length0_re;
	if (videosoc_csrbank1_sram_reader_ev_enable0_re) begin
		ethmac_reader_eventmanager_storage_full <= videosoc_csrbank1_sram_reader_ev_enable0_r;
	end
	ethmac_reader_eventmanager_re <= videosoc_csrbank1_sram_reader_ev_enable0_re;
	videosoc_interface2_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank2_sel) begin
		case (videosoc_interface2_bank_bus_adr[1:0])
			1'd0: begin
				videosoc_interface2_bank_bus_dat_r <= videosoc_csrbank2_crg_reset0_w;
			end
			1'd1: begin
				videosoc_interface2_bank_bus_dat_r <= videosoc_csrbank2_mdio_w0_w;
			end
			2'd2: begin
				videosoc_interface2_bank_bus_dat_r <= videosoc_csrbank2_mdio_r_w;
			end
		endcase
	end
	if (videosoc_csrbank2_crg_reset0_re) begin
		ethphy_reset_storage_full <= videosoc_csrbank2_crg_reset0_r;
	end
	ethphy_reset_re <= videosoc_csrbank2_crg_reset0_re;
	if (videosoc_csrbank2_mdio_w0_re) begin
		ethphy_storage_full[2:0] <= videosoc_csrbank2_mdio_w0_r;
	end
	ethphy_re <= videosoc_csrbank2_mdio_w0_re;
	videosoc_sram0_sel_r <= videosoc_sram0_sel;
	videosoc_interface3_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank3_sel) begin
		case (videosoc_interface3_bank_bus_adr[5:0])
			1'd0: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_edid_hpd_notif_w;
			end
			1'd1: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_edid_hpd_en0_w;
			end
			2'd2: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_mmcm_reset0_w;
			end
			2'd3: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_locked_w;
			end
			3'd4: begin
				videosoc_interface3_bank_bus_dat_r <= mmcm_read_w;
			end
			3'd5: begin
				videosoc_interface3_bank_bus_dat_r <= mmcm_write_w;
			end
			3'd6: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_mmcm_drdy_w;
			end
			3'd7: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_mmcm_adr0_w;
			end
			4'd8: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_mmcm_dat_w1_w;
			end
			4'd9: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_mmcm_dat_w0_w;
			end
			4'd10: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_mmcm_dat_r1_w;
			end
			4'd11: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_clocking_mmcm_dat_r0_w;
			end
			4'd12: begin
				videosoc_interface3_bank_bus_dat_r <= s7datacapture0_dly_ctl_w;
			end
			4'd13: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data0_cap_phase_w;
			end
			4'd14: begin
				videosoc_interface3_bank_bus_dat_r <= s7datacapture0_phase_reset_w;
			end
			4'd15: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data0_charsync_char_synced_w;
			end
			5'd16: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data0_charsync_ctl_pos_w;
			end
			5'd17: begin
				videosoc_interface3_bank_bus_dat_r <= wer0_update_w;
			end
			5'd18: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data0_wer_value2_w;
			end
			5'd19: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data0_wer_value1_w;
			end
			5'd20: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data0_wer_value0_w;
			end
			5'd21: begin
				videosoc_interface3_bank_bus_dat_r <= s7datacapture1_dly_ctl_w;
			end
			5'd22: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data1_cap_phase_w;
			end
			5'd23: begin
				videosoc_interface3_bank_bus_dat_r <= s7datacapture1_phase_reset_w;
			end
			5'd24: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data1_charsync_char_synced_w;
			end
			5'd25: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data1_charsync_ctl_pos_w;
			end
			5'd26: begin
				videosoc_interface3_bank_bus_dat_r <= wer1_update_w;
			end
			5'd27: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data1_wer_value2_w;
			end
			5'd28: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data1_wer_value1_w;
			end
			5'd29: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data1_wer_value0_w;
			end
			5'd30: begin
				videosoc_interface3_bank_bus_dat_r <= s7datacapture2_dly_ctl_w;
			end
			5'd31: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data2_cap_phase_w;
			end
			6'd32: begin
				videosoc_interface3_bank_bus_dat_r <= s7datacapture2_phase_reset_w;
			end
			6'd33: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data2_charsync_char_synced_w;
			end
			6'd34: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data2_charsync_ctl_pos_w;
			end
			6'd35: begin
				videosoc_interface3_bank_bus_dat_r <= wer2_update_w;
			end
			6'd36: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data2_wer_value2_w;
			end
			6'd37: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data2_wer_value1_w;
			end
			6'd38: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_data2_wer_value0_w;
			end
			6'd39: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_chansync_channels_synced_w;
			end
			6'd40: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_resdetection_hres1_w;
			end
			6'd41: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_resdetection_hres0_w;
			end
			6'd42: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_resdetection_vres1_w;
			end
			6'd43: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_resdetection_vres0_w;
			end
			6'd44: begin
				videosoc_interface3_bank_bus_dat_r <= frame_overflow_w;
			end
			6'd45: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_frame_size3_w;
			end
			6'd46: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_frame_size2_w;
			end
			6'd47: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_frame_size1_w;
			end
			6'd48: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_frame_size0_w;
			end
			6'd49: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot0_status0_w;
			end
			6'd50: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot0_address3_w;
			end
			6'd51: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot0_address2_w;
			end
			6'd52: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot0_address1_w;
			end
			6'd53: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot0_address0_w;
			end
			6'd54: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot1_status0_w;
			end
			6'd55: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot1_address3_w;
			end
			6'd56: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot1_address2_w;
			end
			6'd57: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot1_address1_w;
			end
			6'd58: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_slot1_address0_w;
			end
			6'd59: begin
				videosoc_interface3_bank_bus_dat_r <= dma_slot_array_status_w;
			end
			6'd60: begin
				videosoc_interface3_bank_bus_dat_r <= dma_slot_array_pending_w;
			end
			6'd61: begin
				videosoc_interface3_bank_bus_dat_r <= videosoc_csrbank3_dma_ev_enable0_w;
			end
		endcase
	end
	if (videosoc_csrbank3_edid_hpd_en0_re) begin
		edid_storage_full <= videosoc_csrbank3_edid_hpd_en0_r;
	end
	edid_re <= videosoc_csrbank3_edid_hpd_en0_re;
	if (videosoc_csrbank3_clocking_mmcm_reset0_re) begin
		mmcm_reset_storage_full <= videosoc_csrbank3_clocking_mmcm_reset0_r;
	end
	mmcm_reset_re <= videosoc_csrbank3_clocking_mmcm_reset0_re;
	if (videosoc_csrbank3_clocking_mmcm_adr0_re) begin
		mmcm_adr_storage_full[6:0] <= videosoc_csrbank3_clocking_mmcm_adr0_r;
	end
	mmcm_adr_re <= videosoc_csrbank3_clocking_mmcm_adr0_re;
	if (videosoc_csrbank3_clocking_mmcm_dat_w1_re) begin
		mmcm_dat_w_storage_full[15:8] <= videosoc_csrbank3_clocking_mmcm_dat_w1_r;
	end
	if (videosoc_csrbank3_clocking_mmcm_dat_w0_re) begin
		mmcm_dat_w_storage_full[7:0] <= videosoc_csrbank3_clocking_mmcm_dat_w0_r;
	end
	mmcm_dat_w_re <= videosoc_csrbank3_clocking_mmcm_dat_w0_re;
	if (videosoc_csrbank3_dma_frame_size3_re) begin
		dma_frame_size_storage_full[28:24] <= videosoc_csrbank3_dma_frame_size3_r;
	end
	if (videosoc_csrbank3_dma_frame_size2_re) begin
		dma_frame_size_storage_full[23:16] <= videosoc_csrbank3_dma_frame_size2_r;
	end
	if (videosoc_csrbank3_dma_frame_size1_re) begin
		dma_frame_size_storage_full[15:8] <= videosoc_csrbank3_dma_frame_size1_r;
	end
	if (videosoc_csrbank3_dma_frame_size0_re) begin
		dma_frame_size_storage_full[7:0] <= videosoc_csrbank3_dma_frame_size0_r;
	end
	dma_frame_size_re <= videosoc_csrbank3_dma_frame_size0_re;
	if (dma_slot_array_slot0_status_we) begin
		dma_slot_array_slot0_status_storage_full <= (dma_slot_array_slot0_status_dat_w <<< 1'd0);
	end
	if (videosoc_csrbank3_dma_slot0_status0_re) begin
		dma_slot_array_slot0_status_storage_full[1:0] <= videosoc_csrbank3_dma_slot0_status0_r;
	end
	dma_slot_array_slot0_status_re <= videosoc_csrbank3_dma_slot0_status0_re;
	if (dma_slot_array_slot0_address_we) begin
		dma_slot_array_slot0_address_storage_full <= (dma_slot_array_slot0_address_dat_w <<< 3'd4);
	end
	if (videosoc_csrbank3_dma_slot0_address3_re) begin
		dma_slot_array_slot0_address_storage_full[28:24] <= videosoc_csrbank3_dma_slot0_address3_r;
	end
	if (videosoc_csrbank3_dma_slot0_address2_re) begin
		dma_slot_array_slot0_address_storage_full[23:16] <= videosoc_csrbank3_dma_slot0_address2_r;
	end
	if (videosoc_csrbank3_dma_slot0_address1_re) begin
		dma_slot_array_slot0_address_storage_full[15:8] <= videosoc_csrbank3_dma_slot0_address1_r;
	end
	if (videosoc_csrbank3_dma_slot0_address0_re) begin
		dma_slot_array_slot0_address_storage_full[7:0] <= videosoc_csrbank3_dma_slot0_address0_r;
	end
	dma_slot_array_slot0_address_re <= videosoc_csrbank3_dma_slot0_address0_re;
	if (dma_slot_array_slot1_status_we) begin
		dma_slot_array_slot1_status_storage_full <= (dma_slot_array_slot1_status_dat_w <<< 1'd0);
	end
	if (videosoc_csrbank3_dma_slot1_status0_re) begin
		dma_slot_array_slot1_status_storage_full[1:0] <= videosoc_csrbank3_dma_slot1_status0_r;
	end
	dma_slot_array_slot1_status_re <= videosoc_csrbank3_dma_slot1_status0_re;
	if (dma_slot_array_slot1_address_we) begin
		dma_slot_array_slot1_address_storage_full <= (dma_slot_array_slot1_address_dat_w <<< 3'd4);
	end
	if (videosoc_csrbank3_dma_slot1_address3_re) begin
		dma_slot_array_slot1_address_storage_full[28:24] <= videosoc_csrbank3_dma_slot1_address3_r;
	end
	if (videosoc_csrbank3_dma_slot1_address2_re) begin
		dma_slot_array_slot1_address_storage_full[23:16] <= videosoc_csrbank3_dma_slot1_address2_r;
	end
	if (videosoc_csrbank3_dma_slot1_address1_re) begin
		dma_slot_array_slot1_address_storage_full[15:8] <= videosoc_csrbank3_dma_slot1_address1_r;
	end
	if (videosoc_csrbank3_dma_slot1_address0_re) begin
		dma_slot_array_slot1_address_storage_full[7:0] <= videosoc_csrbank3_dma_slot1_address0_r;
	end
	dma_slot_array_slot1_address_re <= videosoc_csrbank3_dma_slot1_address0_re;
	if (videosoc_csrbank3_dma_ev_enable0_re) begin
		dma_slot_array_storage_full[1:0] <= videosoc_csrbank3_dma_ev_enable0_r;
	end
	dma_slot_array_re <= videosoc_csrbank3_dma_ev_enable0_re;
	videosoc_interface4_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank4_sel) begin
		case (videosoc_interface4_bank_bus_adr[1:0])
			1'd0: begin
				videosoc_interface4_bank_bus_dat_r <= videosoc_csrbank4_value3_w;
			end
			1'd1: begin
				videosoc_interface4_bank_bus_dat_r <= videosoc_csrbank4_value2_w;
			end
			2'd2: begin
				videosoc_interface4_bank_bus_dat_r <= videosoc_csrbank4_value1_w;
			end
			2'd3: begin
				videosoc_interface4_bank_bus_dat_r <= videosoc_csrbank4_value0_w;
			end
		endcase
	end
	videosoc_interface5_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank5_sel) begin
		case (videosoc_interface5_bank_bus_adr[5:0])
			1'd0: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_underflow_enable0_w;
			end
			1'd1: begin
				videosoc_interface5_bank_bus_dat_r <= hdmi_out0_core_underflow_update_underflow_update_w;
			end
			2'd2: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_underflow_counter3_w;
			end
			2'd3: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_underflow_counter2_w;
			end
			3'd4: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_underflow_counter1_w;
			end
			3'd5: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_underflow_counter0_w;
			end
			3'd6: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_enable0_w;
			end
			3'd7: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hres1_w;
			end
			4'd8: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hres0_w;
			end
			4'd9: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hsync_start1_w;
			end
			4'd10: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hsync_start0_w;
			end
			4'd11: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hsync_end1_w;
			end
			4'd12: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hsync_end0_w;
			end
			4'd13: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hscan1_w;
			end
			4'd14: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_hscan0_w;
			end
			4'd15: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vres1_w;
			end
			5'd16: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vres0_w;
			end
			5'd17: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vsync_start1_w;
			end
			5'd18: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vsync_start0_w;
			end
			5'd19: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vsync_end1_w;
			end
			5'd20: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vsync_end0_w;
			end
			5'd21: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vscan1_w;
			end
			5'd22: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_vscan0_w;
			end
			5'd23: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_base3_w;
			end
			5'd24: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_base2_w;
			end
			5'd25: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_base1_w;
			end
			5'd26: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_base0_w;
			end
			5'd27: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_length3_w;
			end
			5'd28: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_length2_w;
			end
			5'd29: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_length1_w;
			end
			5'd30: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_core_initiator_length0_w;
			end
			5'd31: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_driver_clocking_mmcm_reset0_w;
			end
			6'd32: begin
				videosoc_interface5_bank_bus_dat_r <= hdmi_out0_driver_s7hdmioutclocking_mmcm_read_w;
			end
			6'd33: begin
				videosoc_interface5_bank_bus_dat_r <= hdmi_out0_driver_s7hdmioutclocking_mmcm_write_w;
			end
			6'd34: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_driver_clocking_mmcm_drdy_w;
			end
			6'd35: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_driver_clocking_mmcm_adr0_w;
			end
			6'd36: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_driver_clocking_mmcm_dat_w1_w;
			end
			6'd37: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_driver_clocking_mmcm_dat_w0_w;
			end
			6'd38: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_driver_clocking_mmcm_dat_r1_w;
			end
			6'd39: begin
				videosoc_interface5_bank_bus_dat_r <= videosoc_csrbank5_driver_clocking_mmcm_dat_r0_w;
			end
		endcase
	end
	if (videosoc_csrbank5_core_underflow_enable0_re) begin
		hdmi_out0_core_underflow_enable_storage_full <= videosoc_csrbank5_core_underflow_enable0_r;
	end
	hdmi_out0_core_underflow_enable_re <= videosoc_csrbank5_core_underflow_enable0_re;
	if (videosoc_csrbank5_core_initiator_enable0_re) begin
		hdmi_out0_core_initiator_enable_storage_full <= videosoc_csrbank5_core_initiator_enable0_r;
	end
	hdmi_out0_core_initiator_enable_re <= videosoc_csrbank5_core_initiator_enable0_re;
	if (videosoc_csrbank5_core_initiator_hres1_re) begin
		videosoc_csrbank5_core_initiator_hres_backstore[3:0] <= videosoc_csrbank5_core_initiator_hres1_r;
	end
	if (videosoc_csrbank5_core_initiator_hres0_re) begin
		hdmi_out0_core_initiator_csrstorage0_storage_full <= {videosoc_csrbank5_core_initiator_hres_backstore, videosoc_csrbank5_core_initiator_hres0_r};
	end
	hdmi_out0_core_initiator_csrstorage0_re <= videosoc_csrbank5_core_initiator_hres0_re;
	if (videosoc_csrbank5_core_initiator_hsync_start1_re) begin
		videosoc_csrbank5_core_initiator_hsync_start_backstore[3:0] <= videosoc_csrbank5_core_initiator_hsync_start1_r;
	end
	if (videosoc_csrbank5_core_initiator_hsync_start0_re) begin
		hdmi_out0_core_initiator_csrstorage1_storage_full <= {videosoc_csrbank5_core_initiator_hsync_start_backstore, videosoc_csrbank5_core_initiator_hsync_start0_r};
	end
	hdmi_out0_core_initiator_csrstorage1_re <= videosoc_csrbank5_core_initiator_hsync_start0_re;
	if (videosoc_csrbank5_core_initiator_hsync_end1_re) begin
		videosoc_csrbank5_core_initiator_hsync_end_backstore[3:0] <= videosoc_csrbank5_core_initiator_hsync_end1_r;
	end
	if (videosoc_csrbank5_core_initiator_hsync_end0_re) begin
		hdmi_out0_core_initiator_csrstorage2_storage_full <= {videosoc_csrbank5_core_initiator_hsync_end_backstore, videosoc_csrbank5_core_initiator_hsync_end0_r};
	end
	hdmi_out0_core_initiator_csrstorage2_re <= videosoc_csrbank5_core_initiator_hsync_end0_re;
	if (videosoc_csrbank5_core_initiator_hscan1_re) begin
		videosoc_csrbank5_core_initiator_hscan_backstore[3:0] <= videosoc_csrbank5_core_initiator_hscan1_r;
	end
	if (videosoc_csrbank5_core_initiator_hscan0_re) begin
		hdmi_out0_core_initiator_csrstorage3_storage_full <= {videosoc_csrbank5_core_initiator_hscan_backstore, videosoc_csrbank5_core_initiator_hscan0_r};
	end
	hdmi_out0_core_initiator_csrstorage3_re <= videosoc_csrbank5_core_initiator_hscan0_re;
	if (videosoc_csrbank5_core_initiator_vres1_re) begin
		videosoc_csrbank5_core_initiator_vres_backstore[3:0] <= videosoc_csrbank5_core_initiator_vres1_r;
	end
	if (videosoc_csrbank5_core_initiator_vres0_re) begin
		hdmi_out0_core_initiator_csrstorage4_storage_full <= {videosoc_csrbank5_core_initiator_vres_backstore, videosoc_csrbank5_core_initiator_vres0_r};
	end
	hdmi_out0_core_initiator_csrstorage4_re <= videosoc_csrbank5_core_initiator_vres0_re;
	if (videosoc_csrbank5_core_initiator_vsync_start1_re) begin
		videosoc_csrbank5_core_initiator_vsync_start_backstore[3:0] <= videosoc_csrbank5_core_initiator_vsync_start1_r;
	end
	if (videosoc_csrbank5_core_initiator_vsync_start0_re) begin
		hdmi_out0_core_initiator_csrstorage5_storage_full <= {videosoc_csrbank5_core_initiator_vsync_start_backstore, videosoc_csrbank5_core_initiator_vsync_start0_r};
	end
	hdmi_out0_core_initiator_csrstorage5_re <= videosoc_csrbank5_core_initiator_vsync_start0_re;
	if (videosoc_csrbank5_core_initiator_vsync_end1_re) begin
		videosoc_csrbank5_core_initiator_vsync_end_backstore[3:0] <= videosoc_csrbank5_core_initiator_vsync_end1_r;
	end
	if (videosoc_csrbank5_core_initiator_vsync_end0_re) begin
		hdmi_out0_core_initiator_csrstorage6_storage_full <= {videosoc_csrbank5_core_initiator_vsync_end_backstore, videosoc_csrbank5_core_initiator_vsync_end0_r};
	end
	hdmi_out0_core_initiator_csrstorage6_re <= videosoc_csrbank5_core_initiator_vsync_end0_re;
	if (videosoc_csrbank5_core_initiator_vscan1_re) begin
		videosoc_csrbank5_core_initiator_vscan_backstore[3:0] <= videosoc_csrbank5_core_initiator_vscan1_r;
	end
	if (videosoc_csrbank5_core_initiator_vscan0_re) begin
		hdmi_out0_core_initiator_csrstorage7_storage_full <= {videosoc_csrbank5_core_initiator_vscan_backstore, videosoc_csrbank5_core_initiator_vscan0_r};
	end
	hdmi_out0_core_initiator_csrstorage7_re <= videosoc_csrbank5_core_initiator_vscan0_re;
	if (videosoc_csrbank5_core_initiator_base3_re) begin
		videosoc_csrbank5_core_initiator_base_backstore[23:16] <= videosoc_csrbank5_core_initiator_base3_r;
	end
	if (videosoc_csrbank5_core_initiator_base2_re) begin
		videosoc_csrbank5_core_initiator_base_backstore[15:8] <= videosoc_csrbank5_core_initiator_base2_r;
	end
	if (videosoc_csrbank5_core_initiator_base1_re) begin
		videosoc_csrbank5_core_initiator_base_backstore[7:0] <= videosoc_csrbank5_core_initiator_base1_r;
	end
	if (videosoc_csrbank5_core_initiator_base0_re) begin
		hdmi_out0_core_initiator_csrstorage8_storage_full <= {videosoc_csrbank5_core_initiator_base_backstore, videosoc_csrbank5_core_initiator_base0_r};
	end
	hdmi_out0_core_initiator_csrstorage8_re <= videosoc_csrbank5_core_initiator_base0_re;
	if (videosoc_csrbank5_core_initiator_length3_re) begin
		videosoc_csrbank5_core_initiator_length_backstore[23:16] <= videosoc_csrbank5_core_initiator_length3_r;
	end
	if (videosoc_csrbank5_core_initiator_length2_re) begin
		videosoc_csrbank5_core_initiator_length_backstore[15:8] <= videosoc_csrbank5_core_initiator_length2_r;
	end
	if (videosoc_csrbank5_core_initiator_length1_re) begin
		videosoc_csrbank5_core_initiator_length_backstore[7:0] <= videosoc_csrbank5_core_initiator_length1_r;
	end
	if (videosoc_csrbank5_core_initiator_length0_re) begin
		hdmi_out0_core_initiator_csrstorage9_storage_full <= {videosoc_csrbank5_core_initiator_length_backstore, videosoc_csrbank5_core_initiator_length0_r};
	end
	hdmi_out0_core_initiator_csrstorage9_re <= videosoc_csrbank5_core_initiator_length0_re;
	if (videosoc_csrbank5_driver_clocking_mmcm_reset0_re) begin
		hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full <= videosoc_csrbank5_driver_clocking_mmcm_reset0_r;
	end
	hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_re <= videosoc_csrbank5_driver_clocking_mmcm_reset0_re;
	if (videosoc_csrbank5_driver_clocking_mmcm_adr0_re) begin
		hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full[6:0] <= videosoc_csrbank5_driver_clocking_mmcm_adr0_r;
	end
	hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_re <= videosoc_csrbank5_driver_clocking_mmcm_adr0_re;
	if (videosoc_csrbank5_driver_clocking_mmcm_dat_w1_re) begin
		hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[15:8] <= videosoc_csrbank5_driver_clocking_mmcm_dat_w1_r;
	end
	if (videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re) begin
		hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[7:0] <= videosoc_csrbank5_driver_clocking_mmcm_dat_w0_r;
	end
	hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_re <= videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re;
	videosoc_sram1_sel_r <= videosoc_sram1_sel;
	videosoc_interface6_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank6_sel) begin
		case (videosoc_interface6_bank_bus_adr[5:0])
			1'd0: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id7_w;
			end
			1'd1: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id6_w;
			end
			2'd2: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id5_w;
			end
			2'd3: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id4_w;
			end
			3'd4: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id3_w;
			end
			3'd5: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id2_w;
			end
			3'd6: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id1_w;
			end
			3'd7: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_dna_id0_w;
			end
			4'd8: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit19_w;
			end
			4'd9: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit18_w;
			end
			4'd10: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit17_w;
			end
			4'd11: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit16_w;
			end
			4'd12: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit15_w;
			end
			4'd13: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit14_w;
			end
			4'd14: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit13_w;
			end
			4'd15: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit12_w;
			end
			5'd16: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit11_w;
			end
			5'd17: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit10_w;
			end
			5'd18: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit9_w;
			end
			5'd19: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit8_w;
			end
			5'd20: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit7_w;
			end
			5'd21: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit6_w;
			end
			5'd22: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit5_w;
			end
			5'd23: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit4_w;
			end
			5'd24: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit3_w;
			end
			5'd25: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit2_w;
			end
			5'd26: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit1_w;
			end
			5'd27: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_git_commit0_w;
			end
			5'd28: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform7_w;
			end
			5'd29: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform6_w;
			end
			5'd30: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform5_w;
			end
			5'd31: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform4_w;
			end
			6'd32: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform3_w;
			end
			6'd33: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform2_w;
			end
			6'd34: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform1_w;
			end
			6'd35: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_platform0_w;
			end
			6'd36: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target7_w;
			end
			6'd37: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target6_w;
			end
			6'd38: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target5_w;
			end
			6'd39: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target4_w;
			end
			6'd40: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target3_w;
			end
			6'd41: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target2_w;
			end
			6'd42: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target1_w;
			end
			6'd43: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_platform_target0_w;
			end
			6'd44: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_temperature1_w;
			end
			6'd45: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_temperature0_w;
			end
			6'd46: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_vccint1_w;
			end
			6'd47: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_vccint0_w;
			end
			6'd48: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_vccaux1_w;
			end
			6'd49: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_vccaux0_w;
			end
			6'd50: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_vccbram1_w;
			end
			6'd51: begin
				videosoc_interface6_bank_bus_dat_r <= videosoc_csrbank6_xadc_vccbram0_w;
			end
		endcase
	end
	videosoc_interface7_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank7_sel) begin
		case (videosoc_interface7_bank_bus_adr[2:0])
			1'd0: begin
				videosoc_interface7_bank_bus_dat_r <= videosoc_oled_spimaster_ctrl_w;
			end
			1'd1: begin
				videosoc_interface7_bank_bus_dat_r <= videosoc_csrbank7_spi_length0_w;
			end
			2'd2: begin
				videosoc_interface7_bank_bus_dat_r <= videosoc_csrbank7_spi_status_w;
			end
			2'd3: begin
				videosoc_interface7_bank_bus_dat_r <= videosoc_csrbank7_spi_mosi0_w;
			end
			3'd4: begin
				videosoc_interface7_bank_bus_dat_r <= videosoc_csrbank7_gpio_out0_w;
			end
		endcase
	end
	if (videosoc_csrbank7_spi_length0_re) begin
		videosoc_oled_spimaster_length_storage_full[7:0] <= videosoc_csrbank7_spi_length0_r;
	end
	videosoc_oled_spimaster_length_re <= videosoc_csrbank7_spi_length0_re;
	if (videosoc_csrbank7_spi_mosi0_re) begin
		videosoc_oled_spimaster_mosi_storage_full[7:0] <= videosoc_csrbank7_spi_mosi0_r;
	end
	videosoc_oled_spimaster_mosi_re <= videosoc_csrbank7_spi_mosi0_re;
	if (videosoc_csrbank7_gpio_out0_re) begin
		videosoc_oled_storage_full[3:0] <= videosoc_csrbank7_gpio_out0_r;
	end
	videosoc_oled_re <= videosoc_csrbank7_gpio_out0_re;
	videosoc_interface8_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank8_sel) begin
		case (videosoc_interface8_bank_bus_adr[5:0])
			1'd0: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_control0_w;
			end
			1'd1: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_command0_w;
			end
			2'd2: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_sdram_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_address1_w;
			end
			3'd4: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_address0_w;
			end
			3'd5: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_baddress0_w;
			end
			3'd6: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_wrdata3_w;
			end
			3'd7: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_wrdata2_w;
			end
			4'd8: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_wrdata1_w;
			end
			4'd9: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_wrdata0_w;
			end
			4'd10: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_rddata3_w;
			end
			4'd11: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_rddata2_w;
			end
			4'd12: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_rddata1_w;
			end
			4'd13: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi0_rddata0_w;
			end
			4'd14: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_command0_w;
			end
			4'd15: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_sdram_phaseinjector1_command_issue_w;
			end
			5'd16: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_address1_w;
			end
			5'd17: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_address0_w;
			end
			5'd18: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_baddress0_w;
			end
			5'd19: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_wrdata3_w;
			end
			5'd20: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_wrdata2_w;
			end
			5'd21: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_wrdata1_w;
			end
			5'd22: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_wrdata0_w;
			end
			5'd23: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_rddata3_w;
			end
			5'd24: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_rddata2_w;
			end
			5'd25: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_rddata1_w;
			end
			5'd26: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi1_rddata0_w;
			end
			5'd27: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_command0_w;
			end
			5'd28: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_sdram_phaseinjector2_command_issue_w;
			end
			5'd29: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_address1_w;
			end
			5'd30: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_address0_w;
			end
			5'd31: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_baddress0_w;
			end
			6'd32: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_wrdata3_w;
			end
			6'd33: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_wrdata2_w;
			end
			6'd34: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_wrdata1_w;
			end
			6'd35: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_wrdata0_w;
			end
			6'd36: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_rddata3_w;
			end
			6'd37: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_rddata2_w;
			end
			6'd38: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_rddata1_w;
			end
			6'd39: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi2_rddata0_w;
			end
			6'd40: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_command0_w;
			end
			6'd41: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_sdram_phaseinjector3_command_issue_w;
			end
			6'd42: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_address1_w;
			end
			6'd43: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_address0_w;
			end
			6'd44: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_baddress0_w;
			end
			6'd45: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_wrdata3_w;
			end
			6'd46: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_wrdata2_w;
			end
			6'd47: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_wrdata1_w;
			end
			6'd48: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_wrdata0_w;
			end
			6'd49: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_rddata3_w;
			end
			6'd50: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_rddata2_w;
			end
			6'd51: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_rddata1_w;
			end
			6'd52: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_dfii_pi3_rddata0_w;
			end
			6'd53: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_sdram_bandwidth_update_w;
			end
			6'd54: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_controller_bandwidth_nreads2_w;
			end
			6'd55: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_controller_bandwidth_nreads1_w;
			end
			6'd56: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_controller_bandwidth_nreads0_w;
			end
			6'd57: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_controller_bandwidth_nwrites2_w;
			end
			6'd58: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_controller_bandwidth_nwrites1_w;
			end
			6'd59: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_controller_bandwidth_nwrites0_w;
			end
			6'd60: begin
				videosoc_interface8_bank_bus_dat_r <= videosoc_csrbank8_controller_bandwidth_data_width_w;
			end
		endcase
	end
	if (videosoc_csrbank8_dfii_control0_re) begin
		videosoc_sdram_storage_full[3:0] <= videosoc_csrbank8_dfii_control0_r;
	end
	videosoc_sdram_re <= videosoc_csrbank8_dfii_control0_re;
	if (videosoc_csrbank8_dfii_pi0_command0_re) begin
		videosoc_sdram_phaseinjector0_command_storage_full[5:0] <= videosoc_csrbank8_dfii_pi0_command0_r;
	end
	videosoc_sdram_phaseinjector0_command_re <= videosoc_csrbank8_dfii_pi0_command0_re;
	if (videosoc_csrbank8_dfii_pi0_address1_re) begin
		videosoc_sdram_phaseinjector0_address_storage_full[14:8] <= videosoc_csrbank8_dfii_pi0_address1_r;
	end
	if (videosoc_csrbank8_dfii_pi0_address0_re) begin
		videosoc_sdram_phaseinjector0_address_storage_full[7:0] <= videosoc_csrbank8_dfii_pi0_address0_r;
	end
	videosoc_sdram_phaseinjector0_address_re <= videosoc_csrbank8_dfii_pi0_address0_re;
	if (videosoc_csrbank8_dfii_pi0_baddress0_re) begin
		videosoc_sdram_phaseinjector0_baddress_storage_full[2:0] <= videosoc_csrbank8_dfii_pi0_baddress0_r;
	end
	videosoc_sdram_phaseinjector0_baddress_re <= videosoc_csrbank8_dfii_pi0_baddress0_re;
	if (videosoc_csrbank8_dfii_pi0_wrdata3_re) begin
		videosoc_sdram_phaseinjector0_wrdata_storage_full[31:24] <= videosoc_csrbank8_dfii_pi0_wrdata3_r;
	end
	if (videosoc_csrbank8_dfii_pi0_wrdata2_re) begin
		videosoc_sdram_phaseinjector0_wrdata_storage_full[23:16] <= videosoc_csrbank8_dfii_pi0_wrdata2_r;
	end
	if (videosoc_csrbank8_dfii_pi0_wrdata1_re) begin
		videosoc_sdram_phaseinjector0_wrdata_storage_full[15:8] <= videosoc_csrbank8_dfii_pi0_wrdata1_r;
	end
	if (videosoc_csrbank8_dfii_pi0_wrdata0_re) begin
		videosoc_sdram_phaseinjector0_wrdata_storage_full[7:0] <= videosoc_csrbank8_dfii_pi0_wrdata0_r;
	end
	videosoc_sdram_phaseinjector0_wrdata_re <= videosoc_csrbank8_dfii_pi0_wrdata0_re;
	if (videosoc_csrbank8_dfii_pi1_command0_re) begin
		videosoc_sdram_phaseinjector1_command_storage_full[5:0] <= videosoc_csrbank8_dfii_pi1_command0_r;
	end
	videosoc_sdram_phaseinjector1_command_re <= videosoc_csrbank8_dfii_pi1_command0_re;
	if (videosoc_csrbank8_dfii_pi1_address1_re) begin
		videosoc_sdram_phaseinjector1_address_storage_full[14:8] <= videosoc_csrbank8_dfii_pi1_address1_r;
	end
	if (videosoc_csrbank8_dfii_pi1_address0_re) begin
		videosoc_sdram_phaseinjector1_address_storage_full[7:0] <= videosoc_csrbank8_dfii_pi1_address0_r;
	end
	videosoc_sdram_phaseinjector1_address_re <= videosoc_csrbank8_dfii_pi1_address0_re;
	if (videosoc_csrbank8_dfii_pi1_baddress0_re) begin
		videosoc_sdram_phaseinjector1_baddress_storage_full[2:0] <= videosoc_csrbank8_dfii_pi1_baddress0_r;
	end
	videosoc_sdram_phaseinjector1_baddress_re <= videosoc_csrbank8_dfii_pi1_baddress0_re;
	if (videosoc_csrbank8_dfii_pi1_wrdata3_re) begin
		videosoc_sdram_phaseinjector1_wrdata_storage_full[31:24] <= videosoc_csrbank8_dfii_pi1_wrdata3_r;
	end
	if (videosoc_csrbank8_dfii_pi1_wrdata2_re) begin
		videosoc_sdram_phaseinjector1_wrdata_storage_full[23:16] <= videosoc_csrbank8_dfii_pi1_wrdata2_r;
	end
	if (videosoc_csrbank8_dfii_pi1_wrdata1_re) begin
		videosoc_sdram_phaseinjector1_wrdata_storage_full[15:8] <= videosoc_csrbank8_dfii_pi1_wrdata1_r;
	end
	if (videosoc_csrbank8_dfii_pi1_wrdata0_re) begin
		videosoc_sdram_phaseinjector1_wrdata_storage_full[7:0] <= videosoc_csrbank8_dfii_pi1_wrdata0_r;
	end
	videosoc_sdram_phaseinjector1_wrdata_re <= videosoc_csrbank8_dfii_pi1_wrdata0_re;
	if (videosoc_csrbank8_dfii_pi2_command0_re) begin
		videosoc_sdram_phaseinjector2_command_storage_full[5:0] <= videosoc_csrbank8_dfii_pi2_command0_r;
	end
	videosoc_sdram_phaseinjector2_command_re <= videosoc_csrbank8_dfii_pi2_command0_re;
	if (videosoc_csrbank8_dfii_pi2_address1_re) begin
		videosoc_sdram_phaseinjector2_address_storage_full[14:8] <= videosoc_csrbank8_dfii_pi2_address1_r;
	end
	if (videosoc_csrbank8_dfii_pi2_address0_re) begin
		videosoc_sdram_phaseinjector2_address_storage_full[7:0] <= videosoc_csrbank8_dfii_pi2_address0_r;
	end
	videosoc_sdram_phaseinjector2_address_re <= videosoc_csrbank8_dfii_pi2_address0_re;
	if (videosoc_csrbank8_dfii_pi2_baddress0_re) begin
		videosoc_sdram_phaseinjector2_baddress_storage_full[2:0] <= videosoc_csrbank8_dfii_pi2_baddress0_r;
	end
	videosoc_sdram_phaseinjector2_baddress_re <= videosoc_csrbank8_dfii_pi2_baddress0_re;
	if (videosoc_csrbank8_dfii_pi2_wrdata3_re) begin
		videosoc_sdram_phaseinjector2_wrdata_storage_full[31:24] <= videosoc_csrbank8_dfii_pi2_wrdata3_r;
	end
	if (videosoc_csrbank8_dfii_pi2_wrdata2_re) begin
		videosoc_sdram_phaseinjector2_wrdata_storage_full[23:16] <= videosoc_csrbank8_dfii_pi2_wrdata2_r;
	end
	if (videosoc_csrbank8_dfii_pi2_wrdata1_re) begin
		videosoc_sdram_phaseinjector2_wrdata_storage_full[15:8] <= videosoc_csrbank8_dfii_pi2_wrdata1_r;
	end
	if (videosoc_csrbank8_dfii_pi2_wrdata0_re) begin
		videosoc_sdram_phaseinjector2_wrdata_storage_full[7:0] <= videosoc_csrbank8_dfii_pi2_wrdata0_r;
	end
	videosoc_sdram_phaseinjector2_wrdata_re <= videosoc_csrbank8_dfii_pi2_wrdata0_re;
	if (videosoc_csrbank8_dfii_pi3_command0_re) begin
		videosoc_sdram_phaseinjector3_command_storage_full[5:0] <= videosoc_csrbank8_dfii_pi3_command0_r;
	end
	videosoc_sdram_phaseinjector3_command_re <= videosoc_csrbank8_dfii_pi3_command0_re;
	if (videosoc_csrbank8_dfii_pi3_address1_re) begin
		videosoc_sdram_phaseinjector3_address_storage_full[14:8] <= videosoc_csrbank8_dfii_pi3_address1_r;
	end
	if (videosoc_csrbank8_dfii_pi3_address0_re) begin
		videosoc_sdram_phaseinjector3_address_storage_full[7:0] <= videosoc_csrbank8_dfii_pi3_address0_r;
	end
	videosoc_sdram_phaseinjector3_address_re <= videosoc_csrbank8_dfii_pi3_address0_re;
	if (videosoc_csrbank8_dfii_pi3_baddress0_re) begin
		videosoc_sdram_phaseinjector3_baddress_storage_full[2:0] <= videosoc_csrbank8_dfii_pi3_baddress0_r;
	end
	videosoc_sdram_phaseinjector3_baddress_re <= videosoc_csrbank8_dfii_pi3_baddress0_re;
	if (videosoc_csrbank8_dfii_pi3_wrdata3_re) begin
		videosoc_sdram_phaseinjector3_wrdata_storage_full[31:24] <= videosoc_csrbank8_dfii_pi3_wrdata3_r;
	end
	if (videosoc_csrbank8_dfii_pi3_wrdata2_re) begin
		videosoc_sdram_phaseinjector3_wrdata_storage_full[23:16] <= videosoc_csrbank8_dfii_pi3_wrdata2_r;
	end
	if (videosoc_csrbank8_dfii_pi3_wrdata1_re) begin
		videosoc_sdram_phaseinjector3_wrdata_storage_full[15:8] <= videosoc_csrbank8_dfii_pi3_wrdata1_r;
	end
	if (videosoc_csrbank8_dfii_pi3_wrdata0_re) begin
		videosoc_sdram_phaseinjector3_wrdata_storage_full[7:0] <= videosoc_csrbank8_dfii_pi3_wrdata0_r;
	end
	videosoc_sdram_phaseinjector3_wrdata_re <= videosoc_csrbank8_dfii_pi3_wrdata0_re;
	videosoc_interface9_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank9_sel) begin
		case (videosoc_interface9_bank_bus_adr[1:0])
			1'd0: begin
				videosoc_interface9_bank_bus_dat_r <= videosoc_csrbank9_bitbang0_w;
			end
			1'd1: begin
				videosoc_interface9_bank_bus_dat_r <= videosoc_csrbank9_miso_w;
			end
			2'd2: begin
				videosoc_interface9_bank_bus_dat_r <= videosoc_csrbank9_bitbang_en0_w;
			end
		endcase
	end
	if (videosoc_csrbank9_bitbang0_re) begin
		videosoc_bitbang_storage_full[3:0] <= videosoc_csrbank9_bitbang0_r;
	end
	videosoc_bitbang_re <= videosoc_csrbank9_bitbang0_re;
	if (videosoc_csrbank9_bitbang_en0_re) begin
		videosoc_bitbang_en_storage_full <= videosoc_csrbank9_bitbang_en0_r;
	end
	videosoc_bitbang_en_re <= videosoc_csrbank9_bitbang_en0_re;
	videosoc_interface10_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank10_sel) begin
		case (videosoc_interface10_bank_bus_adr[4:0])
			1'd0: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_load3_w;
			end
			1'd1: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_load2_w;
			end
			2'd2: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_load1_w;
			end
			2'd3: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_load0_w;
			end
			3'd4: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_reload3_w;
			end
			3'd5: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_reload2_w;
			end
			3'd6: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_reload1_w;
			end
			3'd7: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_reload0_w;
			end
			4'd8: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_en0_w;
			end
			4'd9: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_videosoc_update_value_w;
			end
			4'd10: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_value3_w;
			end
			4'd11: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_value2_w;
			end
			4'd12: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_value1_w;
			end
			4'd13: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_value0_w;
			end
			4'd14: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_videosoc_eventmanager_status_w;
			end
			4'd15: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_videosoc_eventmanager_pending_w;
			end
			5'd16: begin
				videosoc_interface10_bank_bus_dat_r <= videosoc_csrbank10_ev_enable0_w;
			end
		endcase
	end
	if (videosoc_csrbank10_load3_re) begin
		videosoc_videosoc_load_storage_full[31:24] <= videosoc_csrbank10_load3_r;
	end
	if (videosoc_csrbank10_load2_re) begin
		videosoc_videosoc_load_storage_full[23:16] <= videosoc_csrbank10_load2_r;
	end
	if (videosoc_csrbank10_load1_re) begin
		videosoc_videosoc_load_storage_full[15:8] <= videosoc_csrbank10_load1_r;
	end
	if (videosoc_csrbank10_load0_re) begin
		videosoc_videosoc_load_storage_full[7:0] <= videosoc_csrbank10_load0_r;
	end
	videosoc_videosoc_load_re <= videosoc_csrbank10_load0_re;
	if (videosoc_csrbank10_reload3_re) begin
		videosoc_videosoc_reload_storage_full[31:24] <= videosoc_csrbank10_reload3_r;
	end
	if (videosoc_csrbank10_reload2_re) begin
		videosoc_videosoc_reload_storage_full[23:16] <= videosoc_csrbank10_reload2_r;
	end
	if (videosoc_csrbank10_reload1_re) begin
		videosoc_videosoc_reload_storage_full[15:8] <= videosoc_csrbank10_reload1_r;
	end
	if (videosoc_csrbank10_reload0_re) begin
		videosoc_videosoc_reload_storage_full[7:0] <= videosoc_csrbank10_reload0_r;
	end
	videosoc_videosoc_reload_re <= videosoc_csrbank10_reload0_re;
	if (videosoc_csrbank10_en0_re) begin
		videosoc_videosoc_en_storage_full <= videosoc_csrbank10_en0_r;
	end
	videosoc_videosoc_en_re <= videosoc_csrbank10_en0_re;
	if (videosoc_csrbank10_ev_enable0_re) begin
		videosoc_videosoc_eventmanager_storage_full <= videosoc_csrbank10_ev_enable0_r;
	end
	videosoc_videosoc_eventmanager_re <= videosoc_csrbank10_ev_enable0_re;
	videosoc_interface11_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank11_sel) begin
		case (videosoc_interface11_bank_bus_adr[2:0])
			1'd0: begin
				videosoc_interface11_bank_bus_dat_r <= videosoc_uart_rxtx_w;
			end
			1'd1: begin
				videosoc_interface11_bank_bus_dat_r <= videosoc_csrbank11_txfull_w;
			end
			2'd2: begin
				videosoc_interface11_bank_bus_dat_r <= videosoc_csrbank11_rxempty_w;
			end
			2'd3: begin
				videosoc_interface11_bank_bus_dat_r <= videosoc_uart_status_w;
			end
			3'd4: begin
				videosoc_interface11_bank_bus_dat_r <= videosoc_uart_pending_w;
			end
			3'd5: begin
				videosoc_interface11_bank_bus_dat_r <= videosoc_csrbank11_ev_enable0_w;
			end
		endcase
	end
	if (videosoc_csrbank11_ev_enable0_re) begin
		videosoc_uart_storage_full[1:0] <= videosoc_csrbank11_ev_enable0_r;
	end
	videosoc_uart_re <= videosoc_csrbank11_ev_enable0_re;
	videosoc_interface12_bank_bus_dat_r <= 1'd0;
	if (videosoc_csrbank12_sel) begin
		case (videosoc_interface12_bank_bus_adr[1:0])
			1'd0: begin
				videosoc_interface12_bank_bus_dat_r <= videosoc_csrbank12_tuning_word3_w;
			end
			1'd1: begin
				videosoc_interface12_bank_bus_dat_r <= videosoc_csrbank12_tuning_word2_w;
			end
			2'd2: begin
				videosoc_interface12_bank_bus_dat_r <= videosoc_csrbank12_tuning_word1_w;
			end
			2'd3: begin
				videosoc_interface12_bank_bus_dat_r <= videosoc_csrbank12_tuning_word0_w;
			end
		endcase
	end
	if (videosoc_csrbank12_tuning_word3_re) begin
		videosoc_uart_phy_storage_full[31:24] <= videosoc_csrbank12_tuning_word3_r;
	end
	if (videosoc_csrbank12_tuning_word2_re) begin
		videosoc_uart_phy_storage_full[23:16] <= videosoc_csrbank12_tuning_word2_r;
	end
	if (videosoc_csrbank12_tuning_word1_re) begin
		videosoc_uart_phy_storage_full[15:8] <= videosoc_csrbank12_tuning_word1_r;
	end
	if (videosoc_csrbank12_tuning_word0_re) begin
		videosoc_uart_phy_storage_full[7:0] <= videosoc_csrbank12_tuning_word0_r;
	end
	videosoc_uart_phy_re <= videosoc_csrbank12_tuning_word0_re;
	if (sys_rst) begin
		videosoc_videosoc_rom_bus_ack <= 1'd0;
		videosoc_videosoc_sram_bus_ack <= 1'd0;
		videosoc_videosoc_interface_adr <= 14'd0;
		videosoc_videosoc_interface_we <= 1'd0;
		videosoc_videosoc_interface_dat_w <= 8'd0;
		videosoc_videosoc_bus_wishbone_dat_r <= 32'd0;
		videosoc_videosoc_bus_wishbone_ack <= 1'd0;
		videosoc_videosoc_counter <= 2'd0;
		videosoc_videosoc_load_storage_full <= 32'd0;
		videosoc_videosoc_load_re <= 1'd0;
		videosoc_videosoc_reload_storage_full <= 32'd0;
		videosoc_videosoc_reload_re <= 1'd0;
		videosoc_videosoc_en_storage_full <= 1'd0;
		videosoc_videosoc_en_re <= 1'd0;
		videosoc_videosoc_value_status <= 32'd0;
		videosoc_videosoc_zero_pending <= 1'd0;
		videosoc_videosoc_zero_old_trigger <= 1'd0;
		videosoc_videosoc_eventmanager_storage_full <= 1'd0;
		videosoc_videosoc_eventmanager_re <= 1'd0;
		videosoc_videosoc_value <= 32'd0;
		videosoc_uart_tx_pending <= 1'd0;
		videosoc_uart_tx_old_trigger <= 1'd0;
		videosoc_uart_rx_pending <= 1'd0;
		videosoc_uart_rx_old_trigger <= 1'd0;
		videosoc_uart_storage_full <= 2'd0;
		videosoc_uart_re <= 1'd0;
		videosoc_uart_tx_fifo_level <= 5'd0;
		videosoc_uart_tx_fifo_produce <= 4'd0;
		videosoc_uart_tx_fifo_consume <= 4'd0;
		videosoc_uart_rx_fifo_level <= 5'd0;
		videosoc_uart_rx_fifo_produce <= 4'd0;
		videosoc_uart_rx_fifo_consume <= 4'd0;
		videosoc_bridge_count <= 24'd10000000;
		serial_tx <= 1'd1;
		videosoc_uart_phy_storage_full <= 32'd4947802;
		videosoc_uart_phy_re <= 1'd0;
		videosoc_uart_phy_sink_ready <= 1'd0;
		videosoc_uart_phy_uart_clk_txen <= 1'd0;
		videosoc_uart_phy_phase_accumulator_tx <= 32'd0;
		videosoc_uart_phy_tx_reg <= 8'd0;
		videosoc_uart_phy_tx_bitcount <= 4'd0;
		videosoc_uart_phy_tx_busy <= 1'd0;
		videosoc_uart_phy_source_valid <= 1'd0;
		videosoc_uart_phy_uart_clk_rxen <= 1'd0;
		videosoc_uart_phy_phase_accumulator_rx <= 32'd0;
		videosoc_uart_phy_rx_r <= 1'd0;
		videosoc_uart_phy_rx_reg <= 8'd0;
		videosoc_uart_phy_rx_bitcount <= 4'd0;
		videosoc_uart_phy_rx_busy <= 1'd0;
		videosoc_info_dna_status <= 57'd0;
		videosoc_info_dna_cnt <= 7'd0;
		videosoc_info_temperature_status <= 12'd0;
		videosoc_info_vccint_status <= 12'd0;
		videosoc_info_vccaux_status <= 12'd0;
		videosoc_info_vccbram_status <= 12'd0;
		videosoc_oled_spi_pads_clk <= 1'd0;
		videosoc_oled_spi_pads_mosi <= 1'd0;
		videosoc_oled_spimaster_length_storage_full <= 8'd0;
		videosoc_oled_spimaster_length_re <= 1'd0;
		videosoc_oled_spimaster_mosi_storage_full <= 8'd0;
		videosoc_oled_spimaster_mosi_re <= 1'd0;
		videosoc_oled_spimaster_i <= 4'd0;
		videosoc_oled_spimaster_cnt <= 8'd0;
		videosoc_oled_spimaster_sr_mosi <= 8'd0;
		videosoc_oled_storage_full <= 4'd0;
		videosoc_oled_re <= 1'd0;
		videosoc_ddrphy_storage_full <= 2'd0;
		videosoc_ddrphy_re <= 1'd0;
		videosoc_ddrphy_dfi_p0_rddata_valid <= 1'd0;
		videosoc_ddrphy_dfi_p1_rddata_valid <= 1'd0;
		videosoc_ddrphy_dfi_p2_rddata_valid <= 1'd0;
		videosoc_ddrphy_dfi_p3_rddata_valid <= 1'd0;
		videosoc_ddrphy_oe_dqs <= 1'd0;
		videosoc_ddrphy_oe_dq <= 1'd0;
		videosoc_ddrphy_n_rddata_en0 <= 1'd0;
		videosoc_ddrphy_n_rddata_en1 <= 1'd0;
		videosoc_ddrphy_n_rddata_en2 <= 1'd0;
		videosoc_ddrphy_n_rddata_en3 <= 1'd0;
		videosoc_ddrphy_n_rddata_en4 <= 1'd0;
		videosoc_ddrphy_last_wrdata_en <= 4'd0;
		videosoc_sdram_storage_full <= 4'd0;
		videosoc_sdram_re <= 1'd0;
		videosoc_sdram_phaseinjector0_command_storage_full <= 6'd0;
		videosoc_sdram_phaseinjector0_command_re <= 1'd0;
		videosoc_sdram_phaseinjector0_address_storage_full <= 15'd0;
		videosoc_sdram_phaseinjector0_address_re <= 1'd0;
		videosoc_sdram_phaseinjector0_baddress_storage_full <= 3'd0;
		videosoc_sdram_phaseinjector0_baddress_re <= 1'd0;
		videosoc_sdram_phaseinjector0_wrdata_storage_full <= 32'd0;
		videosoc_sdram_phaseinjector0_wrdata_re <= 1'd0;
		videosoc_sdram_phaseinjector0_status <= 32'd0;
		videosoc_sdram_phaseinjector1_command_storage_full <= 6'd0;
		videosoc_sdram_phaseinjector1_command_re <= 1'd0;
		videosoc_sdram_phaseinjector1_address_storage_full <= 15'd0;
		videosoc_sdram_phaseinjector1_address_re <= 1'd0;
		videosoc_sdram_phaseinjector1_baddress_storage_full <= 3'd0;
		videosoc_sdram_phaseinjector1_baddress_re <= 1'd0;
		videosoc_sdram_phaseinjector1_wrdata_storage_full <= 32'd0;
		videosoc_sdram_phaseinjector1_wrdata_re <= 1'd0;
		videosoc_sdram_phaseinjector1_status <= 32'd0;
		videosoc_sdram_phaseinjector2_command_storage_full <= 6'd0;
		videosoc_sdram_phaseinjector2_command_re <= 1'd0;
		videosoc_sdram_phaseinjector2_address_storage_full <= 15'd0;
		videosoc_sdram_phaseinjector2_address_re <= 1'd0;
		videosoc_sdram_phaseinjector2_baddress_storage_full <= 3'd0;
		videosoc_sdram_phaseinjector2_baddress_re <= 1'd0;
		videosoc_sdram_phaseinjector2_wrdata_storage_full <= 32'd0;
		videosoc_sdram_phaseinjector2_wrdata_re <= 1'd0;
		videosoc_sdram_phaseinjector2_status <= 32'd0;
		videosoc_sdram_phaseinjector3_command_storage_full <= 6'd0;
		videosoc_sdram_phaseinjector3_command_re <= 1'd0;
		videosoc_sdram_phaseinjector3_address_storage_full <= 15'd0;
		videosoc_sdram_phaseinjector3_address_re <= 1'd0;
		videosoc_sdram_phaseinjector3_baddress_storage_full <= 3'd0;
		videosoc_sdram_phaseinjector3_baddress_re <= 1'd0;
		videosoc_sdram_phaseinjector3_wrdata_storage_full <= 32'd0;
		videosoc_sdram_phaseinjector3_wrdata_re <= 1'd0;
		videosoc_sdram_phaseinjector3_status <= 32'd0;
		videosoc_sdram_dfi_p0_cas_n <= 1'd1;
		videosoc_sdram_dfi_p0_ras_n <= 1'd1;
		videosoc_sdram_dfi_p0_we_n <= 1'd1;
		videosoc_sdram_dfi_p0_wrdata_en <= 1'd0;
		videosoc_sdram_dfi_p0_rddata_en <= 1'd0;
		videosoc_sdram_dfi_p1_cas_n <= 1'd1;
		videosoc_sdram_dfi_p1_ras_n <= 1'd1;
		videosoc_sdram_dfi_p1_we_n <= 1'd1;
		videosoc_sdram_dfi_p1_wrdata_en <= 1'd0;
		videosoc_sdram_dfi_p1_rddata_en <= 1'd0;
		videosoc_sdram_dfi_p2_cas_n <= 1'd1;
		videosoc_sdram_dfi_p2_ras_n <= 1'd1;
		videosoc_sdram_dfi_p2_we_n <= 1'd1;
		videosoc_sdram_dfi_p2_wrdata_en <= 1'd0;
		videosoc_sdram_dfi_p2_rddata_en <= 1'd0;
		videosoc_sdram_dfi_p3_cas_n <= 1'd1;
		videosoc_sdram_dfi_p3_ras_n <= 1'd1;
		videosoc_sdram_dfi_p3_we_n <= 1'd1;
		videosoc_sdram_dfi_p3_wrdata_en <= 1'd0;
		videosoc_sdram_dfi_p3_rddata_en <= 1'd0;
		videosoc_sdram_seq_done <= 1'd0;
		videosoc_sdram_counter <= 5'd0;
		videosoc_sdram_count <= 10'd782;
		videosoc_sdram_bankmachine0_level <= 4'd0;
		videosoc_sdram_bankmachine0_produce <= 3'd0;
		videosoc_sdram_bankmachine0_consume <= 3'd0;
		videosoc_sdram_bankmachine0_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine0_count <= 3'd5;
		videosoc_sdram_bankmachine1_level <= 4'd0;
		videosoc_sdram_bankmachine1_produce <= 3'd0;
		videosoc_sdram_bankmachine1_consume <= 3'd0;
		videosoc_sdram_bankmachine1_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine1_count <= 3'd5;
		videosoc_sdram_bankmachine2_level <= 4'd0;
		videosoc_sdram_bankmachine2_produce <= 3'd0;
		videosoc_sdram_bankmachine2_consume <= 3'd0;
		videosoc_sdram_bankmachine2_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine2_count <= 3'd5;
		videosoc_sdram_bankmachine3_level <= 4'd0;
		videosoc_sdram_bankmachine3_produce <= 3'd0;
		videosoc_sdram_bankmachine3_consume <= 3'd0;
		videosoc_sdram_bankmachine3_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine3_count <= 3'd5;
		videosoc_sdram_bankmachine4_level <= 4'd0;
		videosoc_sdram_bankmachine4_produce <= 3'd0;
		videosoc_sdram_bankmachine4_consume <= 3'd0;
		videosoc_sdram_bankmachine4_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine4_count <= 3'd5;
		videosoc_sdram_bankmachine5_level <= 4'd0;
		videosoc_sdram_bankmachine5_produce <= 3'd0;
		videosoc_sdram_bankmachine5_consume <= 3'd0;
		videosoc_sdram_bankmachine5_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine5_count <= 3'd5;
		videosoc_sdram_bankmachine6_level <= 4'd0;
		videosoc_sdram_bankmachine6_produce <= 3'd0;
		videosoc_sdram_bankmachine6_consume <= 3'd0;
		videosoc_sdram_bankmachine6_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine6_count <= 3'd5;
		videosoc_sdram_bankmachine7_level <= 4'd0;
		videosoc_sdram_bankmachine7_produce <= 3'd0;
		videosoc_sdram_bankmachine7_consume <= 3'd0;
		videosoc_sdram_bankmachine7_has_openrow <= 1'd0;
		videosoc_sdram_bankmachine7_count <= 3'd5;
		videosoc_sdram_choose_cmd_grant <= 3'd0;
		videosoc_sdram_choose_req_grant <= 3'd0;
		videosoc_sdram_time0 <= 5'd0;
		videosoc_sdram_time1 <= 4'd0;
		videosoc_sdram_bandwidth_nreads_status <= 24'd0;
		videosoc_sdram_bandwidth_nwrites_status <= 24'd0;
		videosoc_sdram_bandwidth_cmd_valid <= 1'd0;
		videosoc_sdram_bandwidth_cmd_ready <= 1'd0;
		videosoc_sdram_bandwidth_cmd_is_read <= 1'd0;
		videosoc_sdram_bandwidth_cmd_is_write <= 1'd0;
		videosoc_sdram_bandwidth_counter <= 24'd0;
		videosoc_sdram_bandwidth_period <= 1'd0;
		videosoc_sdram_bandwidth_nreads <= 24'd0;
		videosoc_sdram_bandwidth_nwrites <= 24'd0;
		videosoc_sdram_bandwidth_nreads_r <= 24'd0;
		videosoc_sdram_bandwidth_nwrites_r <= 24'd0;
		videosoc_adr_offset_r <= 2'd0;
		videosoc_bus_ack <= 1'd0;
		videosoc_bitbang_storage_full <= 4'd0;
		videosoc_bitbang_re <= 1'd0;
		videosoc_bitbang_en_storage_full <= 1'd0;
		videosoc_bitbang_en_re <= 1'd0;
		videosoc_cs_n <= 1'd1;
		videosoc_clk1 <= 1'd0;
		videosoc_sr <= 32'd0;
		videosoc_i <= 1'd0;
		videosoc_miso <= 1'd0;
		videosoc_counter <= 8'd0;
		ethphy_reset_storage_full <= 1'd0;
		ethphy_reset_re <= 1'd0;
		ethphy_counter <= 9'd0;
		ethphy_storage_full <= 3'd0;
		ethphy_re <= 1'd0;
		ethmac_preamble_errors_status <= 32'd0;
		ethmac_crc_errors_status <= 32'd0;
		ethmac_tx_cdc_graycounter0_q <= 7'd0;
		ethmac_tx_cdc_graycounter0_q_binary <= 7'd0;
		ethmac_rx_cdc_graycounter1_q <= 7'd0;
		ethmac_rx_cdc_graycounter1_q_binary <= 7'd0;
		ethmac_writer_errors_status <= 32'd0;
		ethmac_writer_storage_full <= 1'd0;
		ethmac_writer_re <= 1'd0;
		ethmac_writer_counter <= 32'd0;
		ethmac_writer_slot <= 1'd0;
		ethmac_writer_fifo_level <= 2'd0;
		ethmac_writer_fifo_produce <= 1'd0;
		ethmac_writer_fifo_consume <= 1'd0;
		ethmac_reader_slot_storage_full <= 1'd0;
		ethmac_reader_slot_re <= 1'd0;
		ethmac_reader_length_storage_full <= 11'd0;
		ethmac_reader_length_re <= 1'd0;
		ethmac_reader_done_pending <= 1'd0;
		ethmac_reader_eventmanager_storage_full <= 1'd0;
		ethmac_reader_eventmanager_re <= 1'd0;
		ethmac_reader_fifo_level <= 2'd0;
		ethmac_reader_fifo_produce <= 1'd0;
		ethmac_reader_fifo_consume <= 1'd0;
		ethmac_reader_counter <= 11'd0;
		ethmac_reader_last_d <= 1'd0;
		ethmac_sram0_bus_ack0 <= 1'd0;
		ethmac_sram1_bus_ack0 <= 1'd0;
		ethmac_sram0_bus_ack1 <= 1'd0;
		ethmac_sram1_bus_ack1 <= 1'd0;
		ethmac_slave_sel_r <= 4'd0;
		edid_storage_full <= 1'd0;
		edid_re <= 1'd0;
		edid_sda_i <= 1'd0;
		edid_sda_drv_reg <= 1'd0;
		edid_scl_i <= 1'd0;
		edid_samp_count <= 6'd0;
		edid_samp_carry <= 1'd0;
		edid_scl_r <= 1'd0;
		edid_sda_r <= 1'd0;
		edid_din <= 8'd0;
		edid_counter <= 4'd0;
		edid_is_read <= 1'd0;
		edid_offset_counter <= 7'd0;
		edid_data_bit <= 1'd0;
		edid_data_drv <= 1'd0;
		mmcm_reset_storage_full <= 1'd1;
		mmcm_reset_re <= 1'd0;
		mmcm_drdy_status <= 1'd0;
		mmcm_adr_storage_full <= 7'd0;
		mmcm_adr_re <= 1'd0;
		mmcm_dat_w_storage_full <= 16'd0;
		mmcm_dat_w_re <= 1'd0;
		wer0_status <= 24'd0;
		wer0_wer_counter_sys <= 24'd0;
		wer1_status <= 24'd0;
		wer1_wer_counter_sys <= 24'd0;
		wer2_status <= 24'd0;
		wer2_wer_counter_sys <= 24'd0;
		frame_fifo_graycounter1_q <= 10'd0;
		frame_fifo_graycounter1_q_binary <= 10'd0;
		frame_overflow_mask <= 1'd0;
		dma_frame_size_storage_full <= 29'd0;
		dma_frame_size_re <= 1'd0;
		dma_slot_array_slot0_status_storage_full <= 2'd0;
		dma_slot_array_slot0_status_re <= 1'd0;
		dma_slot_array_slot0_address_storage_full <= 29'd0;
		dma_slot_array_slot0_address_re <= 1'd0;
		dma_slot_array_slot1_status_storage_full <= 2'd0;
		dma_slot_array_slot1_status_re <= 1'd0;
		dma_slot_array_slot1_address_storage_full <= 29'd0;
		dma_slot_array_slot1_address_re <= 1'd0;
		dma_slot_array_storage_full <= 2'd0;
		dma_slot_array_re <= 1'd0;
		dma_slot_array_current_slot <= 1'd0;
		dma_current_address <= 25'd0;
		dma_mwords_remaining <= 25'd0;
		dma_fifo_level <= 5'd0;
		dma_fifo_produce <= 4'd0;
		dma_fifo_consume <= 4'd0;
		hdmi_in0_freq_period_counter <= 32'd0;
		hdmi_in0_freq_sampler_o <= 32'd0;
		hdmi_in0_freq_sampler_counter <= 32'd0;
		hdmi_in0_freq_sampler_i_d <= 6'd0;
		hdmi_out0_dram_port_cmd_fifo_graycounter1_q <= 3'd0;
		hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary <= 3'd0;
		hdmi_out0_dram_port_rdata_fifo_graycounter0_q <= 5'd0;
		hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary <= 5'd0;
		hdmi_out0_core_underflow_enable_storage_full <= 1'd0;
		hdmi_out0_core_underflow_enable_re <= 1'd0;
		hdmi_out0_core_initiator_cdc_graycounter0_q <= 2'd0;
		hdmi_out0_core_initiator_cdc_graycounter0_q_binary <= 2'd0;
		hdmi_out0_core_initiator_enable_storage_full <= 1'd0;
		hdmi_out0_core_initiator_enable_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage0_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage0_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage1_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage1_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage2_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage2_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage3_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage3_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage4_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage4_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage5_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage5_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage6_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage6_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage7_storage_full <= 12'd0;
		hdmi_out0_core_initiator_csrstorage7_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage8_storage_full <= 32'd0;
		hdmi_out0_core_initiator_csrstorage8_re <= 1'd0;
		hdmi_out0_core_initiator_csrstorage9_storage_full <= 32'd0;
		hdmi_out0_core_initiator_csrstorage9_re <= 1'd0;
		hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full <= 1'd0;
		hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_re <= 1'd0;
		hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status <= 1'd0;
		hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full <= 7'd0;
		hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_re <= 1'd0;
		hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full <= 16'd0;
		hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_re <= 1'd0;
		wishbonestreamingbridge_state <= 3'd0;
		oled_state <= 2'd0;
		refresher_state <= 2'd0;
		bankmachine0_state <= 3'd0;
		bankmachine1_state <= 3'd0;
		bankmachine2_state <= 3'd0;
		bankmachine3_state <= 3'd0;
		bankmachine4_state <= 3'd0;
		bankmachine5_state <= 3'd0;
		bankmachine6_state <= 3'd0;
		bankmachine7_state <= 3'd0;
		multiplexer_state <= 4'd0;
		roundrobin0_grant <= 2'd0;
		roundrobin1_grant <= 2'd0;
		roundrobin2_grant <= 2'd0;
		roundrobin3_grant <= 2'd0;
		roundrobin4_grant <= 2'd0;
		roundrobin5_grant <= 2'd0;
		roundrobin6_grant <= 2'd0;
		roundrobin7_grant <= 2'd0;
		new_master_wdata_ready0 <= 1'd0;
		new_master_wdata_ready1 <= 1'd0;
		new_master_wdata_ready2 <= 1'd0;
		new_master_wdata_ready3 <= 1'd0;
		new_master_wdata_ready4 <= 1'd0;
		new_master_wdata_ready5 <= 1'd0;
		new_master_wdata_ready6 <= 1'd0;
		new_master_wdata_ready7 <= 1'd0;
		new_master_wdata_ready8 <= 1'd0;
		new_master_rdata_valid0 <= 1'd0;
		new_master_rdata_valid1 <= 1'd0;
		new_master_rdata_valid2 <= 1'd0;
		new_master_rdata_valid3 <= 1'd0;
		new_master_rdata_valid4 <= 1'd0;
		new_master_rdata_valid5 <= 1'd0;
		new_master_rdata_valid6 <= 1'd0;
		new_master_rdata_valid7 <= 1'd0;
		new_master_rdata_valid8 <= 1'd0;
		new_master_rdata_valid9 <= 1'd0;
		new_master_rdata_valid10 <= 1'd0;
		new_master_rdata_valid11 <= 1'd0;
		new_master_rdata_valid12 <= 1'd0;
		new_master_rdata_valid13 <= 1'd0;
		new_master_rdata_valid14 <= 1'd0;
		new_master_rdata_valid15 <= 1'd0;
		new_master_rdata_valid16 <= 1'd0;
		new_master_rdata_valid17 <= 1'd0;
		new_master_rdata_valid18 <= 1'd0;
		new_master_rdata_valid19 <= 1'd0;
		new_master_rdata_valid20 <= 1'd0;
		fullmemorywe_state <= 3'd0;
		litedramwishbonebridge_state <= 2'd0;
		liteethmacsramwriter_state <= 3'd0;
		liteethmacsramreader_state <= 2'd0;
		edid_state <= 4'd0;
		dma_state <= 2'd0;
		videosoc_grant <= 2'd0;
		videosoc_slave_sel_r <= 6'd0;
		videosoc_interface0_bank_bus_dat_r <= 8'd0;
		videosoc_interface1_bank_bus_dat_r <= 8'd0;
		videosoc_interface2_bank_bus_dat_r <= 8'd0;
		videosoc_sram0_sel_r <= 1'd0;
		videosoc_interface3_bank_bus_dat_r <= 8'd0;
		videosoc_interface4_bank_bus_dat_r <= 8'd0;
		videosoc_interface5_bank_bus_dat_r <= 8'd0;
		videosoc_csrbank5_core_initiator_hres_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_hsync_start_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_hsync_end_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_hscan_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_vres_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_vsync_start_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_vsync_end_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_vscan_backstore <= 4'd0;
		videosoc_csrbank5_core_initiator_base_backstore <= 24'd0;
		videosoc_csrbank5_core_initiator_length_backstore <= 24'd0;
		videosoc_sram1_sel_r <= 1'd0;
		videosoc_interface6_bank_bus_dat_r <= 8'd0;
		videosoc_interface7_bank_bus_dat_r <= 8'd0;
		videosoc_interface8_bank_bus_dat_r <= 8'd0;
		videosoc_interface9_bank_bus_dat_r <= 8'd0;
		videosoc_interface10_bank_bus_dat_r <= 8'd0;
		videosoc_interface11_bank_bus_dat_r <= 8'd0;
		videosoc_interface12_bank_bus_dat_r <= 8'd0;
	end
	xilinxmultiregimpl0_regs0 <= serial_rx;
	xilinxmultiregimpl0_regs1 <= xilinxmultiregimpl0_regs0;
	xilinxmultiregimpl1_regs0 <= ethphy_data_r;
	xilinxmultiregimpl1_regs1 <= xilinxmultiregimpl1_regs0;
	xilinxmultiregimpl2_regs0 <= ethmac_ps_preamble_error_toggle_i;
	xilinxmultiregimpl2_regs1 <= xilinxmultiregimpl2_regs0;
	xilinxmultiregimpl3_regs0 <= ethmac_ps_crc_error_toggle_i;
	xilinxmultiregimpl3_regs1 <= xilinxmultiregimpl3_regs0;
	xilinxmultiregimpl5_regs0 <= ethmac_tx_cdc_graycounter1_q;
	xilinxmultiregimpl5_regs1 <= xilinxmultiregimpl5_regs0;
	xilinxmultiregimpl6_regs0 <= ethmac_rx_cdc_graycounter0_q;
	xilinxmultiregimpl6_regs1 <= xilinxmultiregimpl6_regs0;
	xilinxmultiregimpl8_regs0 <= hdmi_in_scl;
	xilinxmultiregimpl8_regs1 <= xilinxmultiregimpl8_regs0;
	xilinxmultiregimpl9_regs0 <= edid_sda_i_async;
	xilinxmultiregimpl9_regs1 <= xilinxmultiregimpl9_regs0;
	xilinxmultiregimpl10_regs0 <= mmcm_locked;
	xilinxmultiregimpl10_regs1 <= xilinxmultiregimpl10_regs0;
	xilinxmultiregimpl16_regs0 <= {s7datacapture0_too_early, s7datacapture0_too_late};
	xilinxmultiregimpl16_regs1 <= xilinxmultiregimpl16_regs0;
	xilinxmultiregimpl18_regs0 <= charsync0_synced;
	xilinxmultiregimpl18_regs1 <= xilinxmultiregimpl18_regs0;
	xilinxmultiregimpl19_regs0 <= charsync0_word_sel;
	xilinxmultiregimpl19_regs1 <= xilinxmultiregimpl19_regs0;
	xilinxmultiregimpl20_regs0 <= wer0_toggle_i;
	xilinxmultiregimpl20_regs1 <= xilinxmultiregimpl20_regs0;
	xilinxmultiregimpl26_regs0 <= {s7datacapture1_too_early, s7datacapture1_too_late};
	xilinxmultiregimpl26_regs1 <= xilinxmultiregimpl26_regs0;
	xilinxmultiregimpl28_regs0 <= charsync1_synced;
	xilinxmultiregimpl28_regs1 <= xilinxmultiregimpl28_regs0;
	xilinxmultiregimpl29_regs0 <= charsync1_word_sel;
	xilinxmultiregimpl29_regs1 <= xilinxmultiregimpl29_regs0;
	xilinxmultiregimpl30_regs0 <= wer1_toggle_i;
	xilinxmultiregimpl30_regs1 <= xilinxmultiregimpl30_regs0;
	xilinxmultiregimpl36_regs0 <= {s7datacapture2_too_early, s7datacapture2_too_late};
	xilinxmultiregimpl36_regs1 <= xilinxmultiregimpl36_regs0;
	xilinxmultiregimpl38_regs0 <= charsync2_synced;
	xilinxmultiregimpl38_regs1 <= xilinxmultiregimpl38_regs0;
	xilinxmultiregimpl39_regs0 <= charsync2_word_sel;
	xilinxmultiregimpl39_regs1 <= xilinxmultiregimpl39_regs0;
	xilinxmultiregimpl40_regs0 <= wer2_toggle_i;
	xilinxmultiregimpl40_regs1 <= xilinxmultiregimpl40_regs0;
	xilinxmultiregimpl41_regs0 <= chansync_chan_synced;
	xilinxmultiregimpl41_regs1 <= xilinxmultiregimpl41_regs0;
	xilinxmultiregimpl42_regs0 <= resdetection_hcounter_st;
	xilinxmultiregimpl42_regs1 <= xilinxmultiregimpl42_regs0;
	xilinxmultiregimpl43_regs0 <= resdetection_vcounter_st;
	xilinxmultiregimpl43_regs1 <= xilinxmultiregimpl43_regs0;
	xilinxmultiregimpl44_regs0 <= frame_fifo_graycounter0_q;
	xilinxmultiregimpl44_regs1 <= xilinxmultiregimpl44_regs0;
	xilinxmultiregimpl46_regs0 <= frame_pix_overflow;
	xilinxmultiregimpl46_regs1 <= xilinxmultiregimpl46_regs0;
	xilinxmultiregimpl48_regs0 <= frame_overflow_reset_ack_toggle_i;
	xilinxmultiregimpl48_regs1 <= xilinxmultiregimpl48_regs0;
	xilinxmultiregimpl49_regs0 <= hdmi_in0_freq_q;
	xilinxmultiregimpl49_regs1 <= xilinxmultiregimpl49_regs0;
	xilinxmultiregimpl50_regs0 <= hdmi_out0_dram_port_cmd_fifo_graycounter0_q;
	xilinxmultiregimpl50_regs1 <= xilinxmultiregimpl50_regs0;
	xilinxmultiregimpl53_regs0 <= hdmi_out0_dram_port_rdata_fifo_graycounter1_q;
	xilinxmultiregimpl53_regs1 <= xilinxmultiregimpl53_regs0;
	xilinxmultiregimpl55_regs0 <= hdmi_out0_core_initiator_cdc_graycounter1_q;
	xilinxmultiregimpl55_regs1 <= xilinxmultiregimpl55_regs0;
	xilinxmultiregimpl56_regs0 <= hdmi_out0_core_underflow_enable_storage;
	xilinxmultiregimpl56_regs1 <= xilinxmultiregimpl56_regs0;
end

lm32_cpu #(
	.eba_reset(32'h00000000)
) lm32_cpu (
	.D_ACK_I(videosoc_videosoc_dbus_ack),
	.D_DAT_I(videosoc_videosoc_dbus_dat_r),
	.D_ERR_I(videosoc_videosoc_dbus_err),
	.D_RTY_I(1'd0),
	.I_ACK_I(videosoc_videosoc_ibus_ack),
	.I_DAT_I(videosoc_videosoc_ibus_dat_r),
	.I_ERR_I(videosoc_videosoc_ibus_err),
	.I_RTY_I(1'd0),
	.clk_i(sys_clk),
	.interrupt(videosoc_videosoc_interrupt),
	.rst_i(sys_rst),
	.D_ADR_O(videosoc_videosoc_d_adr_o),
	.D_BTE_O(videosoc_videosoc_dbus_bte),
	.D_CTI_O(videosoc_videosoc_dbus_cti),
	.D_CYC_O(videosoc_videosoc_dbus_cyc),
	.D_DAT_O(videosoc_videosoc_dbus_dat_w),
	.D_SEL_O(videosoc_videosoc_dbus_sel),
	.D_STB_O(videosoc_videosoc_dbus_stb),
	.D_WE_O(videosoc_videosoc_dbus_we),
	.I_ADR_O(videosoc_videosoc_i_adr_o),
	.I_BTE_O(videosoc_videosoc_ibus_bte),
	.I_CTI_O(videosoc_videosoc_ibus_cti),
	.I_CYC_O(videosoc_videosoc_ibus_cyc),
	.I_DAT_O(videosoc_videosoc_ibus_dat_w),
	.I_SEL_O(videosoc_videosoc_ibus_sel),
	.I_STB_O(videosoc_videosoc_ibus_stb),
	.I_WE_O(videosoc_videosoc_ibus_we)
);

reg [31:0] mem[0:8191];
reg [31:0] memdat;
always @(posedge sys_clk) begin
	memdat <= mem[videosoc_videosoc_rom_adr];
end

assign videosoc_videosoc_rom_dat_r = memdat;

initial begin
	$readmemh("mem.init", mem);
end

reg [31:0] mem_1[0:8191];
reg [12:0] memadr;
always @(posedge sys_clk) begin
	if (videosoc_videosoc_sram_we[0])
		mem_1[videosoc_videosoc_sram_adr][7:0] <= videosoc_videosoc_sram_dat_w[7:0];
	if (videosoc_videosoc_sram_we[1])
		mem_1[videosoc_videosoc_sram_adr][15:8] <= videosoc_videosoc_sram_dat_w[15:8];
	if (videosoc_videosoc_sram_we[2])
		mem_1[videosoc_videosoc_sram_adr][23:16] <= videosoc_videosoc_sram_dat_w[23:16];
	if (videosoc_videosoc_sram_we[3])
		mem_1[videosoc_videosoc_sram_adr][31:24] <= videosoc_videosoc_sram_dat_w[31:24];
	memadr <= videosoc_videosoc_sram_adr;
end

assign videosoc_videosoc_sram_dat_r = mem_1[memadr];

reg [7:0] mem_2[0:8];
reg [7:0] memdat_1;
always @(posedge sys_clk) begin
	memdat_1 <= mem_2[videosoc_sram1_adr];
end

assign videosoc_sram1_dat_r = memdat_1;

initial begin
	$readmemh("mem_2.init", mem_2);
end

PLLE2_BASE #(
	.CLKFBOUT_MULT(5'd16),
	.CLKIN1_PERIOD(10.0),
	.CLKOUT0_DIVIDE(5'd16),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(3'd4),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(3'd4),
	.CLKOUT2_PHASE(90.0),
	.CLKOUT3_DIVIDE(4'd8),
	.CLKOUT3_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_BASE (
	.CLKFBIN(videosoc_pll_fb),
	.CLKIN1(clk100),
	.CLKFBOUT(videosoc_pll_fb),
	.CLKOUT0(videosoc_pll_sys),
	.CLKOUT1(videosoc_pll_sys4x),
	.CLKOUT2(videosoc_pll_sys4x_dqs),
	.CLKOUT3(videosoc_pll_clk200),
	.LOCKED(videosoc_pll_locked)
);

BUFG BUFG(
	.I(videosoc_pll_sys),
	.O(sys_clk)
);

BUFG BUFG_1(
	.I(videosoc_pll_sys4x),
	.O(sys4x_clk)
);

BUFG BUFG_2(
	.I(videosoc_pll_sys4x_dqs),
	.O(sys4x_dqs_clk)
);

BUFG BUFG_3(
	.I(videosoc_pll_clk200),
	.O(clk200_clk)
);

BUFG BUFG_4(
	.I(clk100),
	.O(clk100_clk)
);

IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(videosoc_ic_reset)
);

reg [9:0] storage[0:15];
reg [3:0] memadr_1;
always @(posedge sys_clk) begin
	if (videosoc_uart_tx_fifo_wrport_we)
		storage[videosoc_uart_tx_fifo_wrport_adr] <= videosoc_uart_tx_fifo_wrport_dat_w;
	memadr_1 <= videosoc_uart_tx_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_uart_tx_fifo_wrport_dat_r = storage[memadr_1];
assign videosoc_uart_tx_fifo_rdport_dat_r = storage[videosoc_uart_tx_fifo_rdport_adr];

reg [9:0] storage_1[0:15];
reg [3:0] memadr_2;
always @(posedge sys_clk) begin
	if (videosoc_uart_rx_fifo_wrport_we)
		storage_1[videosoc_uart_rx_fifo_wrport_adr] <= videosoc_uart_rx_fifo_wrport_dat_w;
	memadr_2 <= videosoc_uart_rx_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_uart_rx_fifo_wrport_dat_r = storage_1[memadr_2];
assign videosoc_uart_rx_fifo_rdport_dat_r = storage_1[videosoc_uart_rx_fifo_rdport_adr];

DNA_PORT DNA_PORT(
	.CLK(videosoc_info_dna_cnt[0]),
	.DIN(videosoc_info_dna_status[56]),
	.READ((videosoc_info_dna_cnt < 2'd2)),
	.SHIFT(1'd1),
	.DOUT(videosoc_info_dna_do)
);

XADC #(
	.INIT_40(16'd36864),
	.INIT_41(14'd12016),
	.INIT_42(11'd1024),
	.INIT_48(15'd18177),
	.INIT_49(4'd15),
	.INIT_4A(15'd18176),
	.INIT_4B(1'd0),
	.INIT_4C(1'd0),
	.INIT_4D(1'd0),
	.INIT_4E(1'd0),
	.INIT_4F(1'd0),
	.INIT_50(16'd46573),
	.INIT_51(15'd22937),
	.INIT_52(16'd41287),
	.INIT_53(16'd56797),
	.INIT_54(16'd43322),
	.INIT_55(15'd20753),
	.INIT_56(16'd37355),
	.INIT_57(16'd44622),
	.INIT_58(15'd22937),
	.INIT_5C(15'd20753)
) XADC (
	.CONVST(1'd0),
	.CONVSTCLK(1'd0),
	.DADDR(videosoc_info_channel),
	.DCLK(sys_clk),
	.DEN(videosoc_info_eoc),
	.DI(1'd0),
	.DWE(1'd0),
	.RESET(sys_rst),
	.VAUXN(1'd0),
	.VAUXP(1'd1),
	.VN(1'd0),
	.VP(1'd1),
	.ALM(videosoc_info_alarm),
	.BUSY(videosoc_info_busy),
	.CHANNEL(videosoc_info_channel),
	.DO(videosoc_info_data),
	.DRDY(videosoc_info_drdy),
	.EOC(videosoc_info_eoc),
	.EOS(videosoc_info_eos),
	.OT(videosoc_info_ot)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(videosoc_ddrphy_sd_clk_se)
);

OBUFDS OBUFDS(
	.I(videosoc_ddrphy_sd_clk_se),
	.O(ddram_clk_p),
	.OB(ddram_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[0]),
	.D2(videosoc_ddrphy_dfi_p0_address[0]),
	.D3(videosoc_ddrphy_dfi_p1_address[0]),
	.D4(videosoc_ddrphy_dfi_p1_address[0]),
	.D5(videosoc_ddrphy_dfi_p2_address[0]),
	.D6(videosoc_ddrphy_dfi_p2_address[0]),
	.D7(videosoc_ddrphy_dfi_p3_address[0]),
	.D8(videosoc_ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[1]),
	.D2(videosoc_ddrphy_dfi_p0_address[1]),
	.D3(videosoc_ddrphy_dfi_p1_address[1]),
	.D4(videosoc_ddrphy_dfi_p1_address[1]),
	.D5(videosoc_ddrphy_dfi_p2_address[1]),
	.D6(videosoc_ddrphy_dfi_p2_address[1]),
	.D7(videosoc_ddrphy_dfi_p3_address[1]),
	.D8(videosoc_ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[2]),
	.D2(videosoc_ddrphy_dfi_p0_address[2]),
	.D3(videosoc_ddrphy_dfi_p1_address[2]),
	.D4(videosoc_ddrphy_dfi_p1_address[2]),
	.D5(videosoc_ddrphy_dfi_p2_address[2]),
	.D6(videosoc_ddrphy_dfi_p2_address[2]),
	.D7(videosoc_ddrphy_dfi_p3_address[2]),
	.D8(videosoc_ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[3]),
	.D2(videosoc_ddrphy_dfi_p0_address[3]),
	.D3(videosoc_ddrphy_dfi_p1_address[3]),
	.D4(videosoc_ddrphy_dfi_p1_address[3]),
	.D5(videosoc_ddrphy_dfi_p2_address[3]),
	.D6(videosoc_ddrphy_dfi_p2_address[3]),
	.D7(videosoc_ddrphy_dfi_p3_address[3]),
	.D8(videosoc_ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[4]),
	.D2(videosoc_ddrphy_dfi_p0_address[4]),
	.D3(videosoc_ddrphy_dfi_p1_address[4]),
	.D4(videosoc_ddrphy_dfi_p1_address[4]),
	.D5(videosoc_ddrphy_dfi_p2_address[4]),
	.D6(videosoc_ddrphy_dfi_p2_address[4]),
	.D7(videosoc_ddrphy_dfi_p3_address[4]),
	.D8(videosoc_ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[5]),
	.D2(videosoc_ddrphy_dfi_p0_address[5]),
	.D3(videosoc_ddrphy_dfi_p1_address[5]),
	.D4(videosoc_ddrphy_dfi_p1_address[5]),
	.D5(videosoc_ddrphy_dfi_p2_address[5]),
	.D6(videosoc_ddrphy_dfi_p2_address[5]),
	.D7(videosoc_ddrphy_dfi_p3_address[5]),
	.D8(videosoc_ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[6]),
	.D2(videosoc_ddrphy_dfi_p0_address[6]),
	.D3(videosoc_ddrphy_dfi_p1_address[6]),
	.D4(videosoc_ddrphy_dfi_p1_address[6]),
	.D5(videosoc_ddrphy_dfi_p2_address[6]),
	.D6(videosoc_ddrphy_dfi_p2_address[6]),
	.D7(videosoc_ddrphy_dfi_p3_address[6]),
	.D8(videosoc_ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[7]),
	.D2(videosoc_ddrphy_dfi_p0_address[7]),
	.D3(videosoc_ddrphy_dfi_p1_address[7]),
	.D4(videosoc_ddrphy_dfi_p1_address[7]),
	.D5(videosoc_ddrphy_dfi_p2_address[7]),
	.D6(videosoc_ddrphy_dfi_p2_address[7]),
	.D7(videosoc_ddrphy_dfi_p3_address[7]),
	.D8(videosoc_ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[8]),
	.D2(videosoc_ddrphy_dfi_p0_address[8]),
	.D3(videosoc_ddrphy_dfi_p1_address[8]),
	.D4(videosoc_ddrphy_dfi_p1_address[8]),
	.D5(videosoc_ddrphy_dfi_p2_address[8]),
	.D6(videosoc_ddrphy_dfi_p2_address[8]),
	.D7(videosoc_ddrphy_dfi_p3_address[8]),
	.D8(videosoc_ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[8])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[9]),
	.D2(videosoc_ddrphy_dfi_p0_address[9]),
	.D3(videosoc_ddrphy_dfi_p1_address[9]),
	.D4(videosoc_ddrphy_dfi_p1_address[9]),
	.D5(videosoc_ddrphy_dfi_p2_address[9]),
	.D6(videosoc_ddrphy_dfi_p2_address[9]),
	.D7(videosoc_ddrphy_dfi_p3_address[9]),
	.D8(videosoc_ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[9])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[10]),
	.D2(videosoc_ddrphy_dfi_p0_address[10]),
	.D3(videosoc_ddrphy_dfi_p1_address[10]),
	.D4(videosoc_ddrphy_dfi_p1_address[10]),
	.D5(videosoc_ddrphy_dfi_p2_address[10]),
	.D6(videosoc_ddrphy_dfi_p2_address[10]),
	.D7(videosoc_ddrphy_dfi_p3_address[10]),
	.D8(videosoc_ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[10])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[11]),
	.D2(videosoc_ddrphy_dfi_p0_address[11]),
	.D3(videosoc_ddrphy_dfi_p1_address[11]),
	.D4(videosoc_ddrphy_dfi_p1_address[11]),
	.D5(videosoc_ddrphy_dfi_p2_address[11]),
	.D6(videosoc_ddrphy_dfi_p2_address[11]),
	.D7(videosoc_ddrphy_dfi_p3_address[11]),
	.D8(videosoc_ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[11])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[12]),
	.D2(videosoc_ddrphy_dfi_p0_address[12]),
	.D3(videosoc_ddrphy_dfi_p1_address[12]),
	.D4(videosoc_ddrphy_dfi_p1_address[12]),
	.D5(videosoc_ddrphy_dfi_p2_address[12]),
	.D6(videosoc_ddrphy_dfi_p2_address[12]),
	.D7(videosoc_ddrphy_dfi_p3_address[12]),
	.D8(videosoc_ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[12])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[13]),
	.D2(videosoc_ddrphy_dfi_p0_address[13]),
	.D3(videosoc_ddrphy_dfi_p1_address[13]),
	.D4(videosoc_ddrphy_dfi_p1_address[13]),
	.D5(videosoc_ddrphy_dfi_p2_address[13]),
	.D6(videosoc_ddrphy_dfi_p2_address[13]),
	.D7(videosoc_ddrphy_dfi_p3_address[13]),
	.D8(videosoc_ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[13])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_address[14]),
	.D2(videosoc_ddrphy_dfi_p0_address[14]),
	.D3(videosoc_ddrphy_dfi_p1_address[14]),
	.D4(videosoc_ddrphy_dfi_p1_address[14]),
	.D5(videosoc_ddrphy_dfi_p2_address[14]),
	.D6(videosoc_ddrphy_dfi_p2_address[14]),
	.D7(videosoc_ddrphy_dfi_p3_address[14]),
	.D8(videosoc_ddrphy_dfi_p3_address[14]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[14])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_bank[0]),
	.D2(videosoc_ddrphy_dfi_p0_bank[0]),
	.D3(videosoc_ddrphy_dfi_p1_bank[0]),
	.D4(videosoc_ddrphy_dfi_p1_bank[0]),
	.D5(videosoc_ddrphy_dfi_p2_bank[0]),
	.D6(videosoc_ddrphy_dfi_p2_bank[0]),
	.D7(videosoc_ddrphy_dfi_p3_bank[0]),
	.D8(videosoc_ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_bank[1]),
	.D2(videosoc_ddrphy_dfi_p0_bank[1]),
	.D3(videosoc_ddrphy_dfi_p1_bank[1]),
	.D4(videosoc_ddrphy_dfi_p1_bank[1]),
	.D5(videosoc_ddrphy_dfi_p2_bank[1]),
	.D6(videosoc_ddrphy_dfi_p2_bank[1]),
	.D7(videosoc_ddrphy_dfi_p3_bank[1]),
	.D8(videosoc_ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_bank[2]),
	.D2(videosoc_ddrphy_dfi_p0_bank[2]),
	.D3(videosoc_ddrphy_dfi_p1_bank[2]),
	.D4(videosoc_ddrphy_dfi_p1_bank[2]),
	.D5(videosoc_ddrphy_dfi_p2_bank[2]),
	.D6(videosoc_ddrphy_dfi_p2_bank[2]),
	.D7(videosoc_ddrphy_dfi_p3_bank[2]),
	.D8(videosoc_ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_ras_n),
	.D2(videosoc_ddrphy_dfi_p0_ras_n),
	.D3(videosoc_ddrphy_dfi_p1_ras_n),
	.D4(videosoc_ddrphy_dfi_p1_ras_n),
	.D5(videosoc_ddrphy_dfi_p2_ras_n),
	.D6(videosoc_ddrphy_dfi_p2_ras_n),
	.D7(videosoc_ddrphy_dfi_p3_ras_n),
	.D8(videosoc_ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_cas_n),
	.D2(videosoc_ddrphy_dfi_p0_cas_n),
	.D3(videosoc_ddrphy_dfi_p1_cas_n),
	.D4(videosoc_ddrphy_dfi_p1_cas_n),
	.D5(videosoc_ddrphy_dfi_p2_cas_n),
	.D6(videosoc_ddrphy_dfi_p2_cas_n),
	.D7(videosoc_ddrphy_dfi_p3_cas_n),
	.D8(videosoc_ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_we_n),
	.D2(videosoc_ddrphy_dfi_p0_we_n),
	.D3(videosoc_ddrphy_dfi_p1_we_n),
	.D4(videosoc_ddrphy_dfi_p1_we_n),
	.D5(videosoc_ddrphy_dfi_p2_we_n),
	.D6(videosoc_ddrphy_dfi_p2_we_n),
	.D7(videosoc_ddrphy_dfi_p3_we_n),
	.D8(videosoc_ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_cke),
	.D2(videosoc_ddrphy_dfi_p0_cke),
	.D3(videosoc_ddrphy_dfi_p1_cke),
	.D4(videosoc_ddrphy_dfi_p1_cke),
	.D5(videosoc_ddrphy_dfi_p2_cke),
	.D6(videosoc_ddrphy_dfi_p2_cke),
	.D7(videosoc_ddrphy_dfi_p3_cke),
	.D8(videosoc_ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_odt),
	.D2(videosoc_ddrphy_dfi_p0_odt),
	.D3(videosoc_ddrphy_dfi_p1_odt),
	.D4(videosoc_ddrphy_dfi_p1_odt),
	.D5(videosoc_ddrphy_dfi_p2_odt),
	.D6(videosoc_ddrphy_dfi_p2_odt),
	.D7(videosoc_ddrphy_dfi_p3_odt),
	.D8(videosoc_ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_reset_n),
	.D2(videosoc_ddrphy_dfi_p0_reset_n),
	.D3(videosoc_ddrphy_dfi_p1_reset_n),
	.D4(videosoc_ddrphy_dfi_p1_reset_n),
	.D5(videosoc_ddrphy_dfi_p2_reset_n),
	.D6(videosoc_ddrphy_dfi_p2_reset_n),
	.D7(videosoc_ddrphy_dfi_p3_reset_n),
	.D8(videosoc_ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata_mask[2]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata_mask[2]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata_mask[2]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata_mask[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dqs_serdes_pattern[0]),
	.D2(videosoc_ddrphy_dqs_serdes_pattern[1]),
	.D3(videosoc_ddrphy_dqs_serdes_pattern[2]),
	.D4(videosoc_ddrphy_dqs_serdes_pattern[3]),
	.D5(videosoc_ddrphy_dqs_serdes_pattern[4]),
	.D6(videosoc_ddrphy_dqs_serdes_pattern[5]),
	.D7(videosoc_ddrphy_dqs_serdes_pattern[6]),
	.D8(videosoc_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dqs0),
	.TQ(videosoc_ddrphy_dqs_t0)
);

OBUFTDS OBUFTDS(
	.I(videosoc_ddrphy_dqs0),
	.T(videosoc_ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata_mask[3]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata_mask[3]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata_mask[3]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata_mask[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dqs_serdes_pattern[0]),
	.D2(videosoc_ddrphy_dqs_serdes_pattern[1]),
	.D3(videosoc_ddrphy_dqs_serdes_pattern[2]),
	.D4(videosoc_ddrphy_dqs_serdes_pattern[3]),
	.D5(videosoc_ddrphy_dqs_serdes_pattern[4]),
	.D6(videosoc_ddrphy_dqs_serdes_pattern[5]),
	.D7(videosoc_ddrphy_dqs_serdes_pattern[6]),
	.D8(videosoc_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dqs1),
	.TQ(videosoc_ddrphy_dqs_t1)
);

OBUFTDS OBUFTDS_1(
	.I(videosoc_ddrphy_dqs1),
	.T(videosoc_ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[0]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[16]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[0]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[16]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[0]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[16]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[0]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[16]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o0),
	.TQ(videosoc_ddrphy_dq_t0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed0),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[16]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[0]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[16]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[0]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[16]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[0]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[16]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed0)
);

IOBUF IOBUF(
	.I(videosoc_ddrphy_dq_o0),
	.T(videosoc_ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(videosoc_ddrphy_dq_i_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[1]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[17]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[1]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[17]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[1]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[17]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[1]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[17]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o1),
	.TQ(videosoc_ddrphy_dq_t1)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed1),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[17]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[1]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[17]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[1]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[17]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[1]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[17]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[1])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed1)
);

IOBUF IOBUF_1(
	.I(videosoc_ddrphy_dq_o1),
	.T(videosoc_ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(videosoc_ddrphy_dq_i_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[2]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[18]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[2]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[18]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[2]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[18]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[2]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[18]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o2),
	.TQ(videosoc_ddrphy_dq_t2)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed2),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[18]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[2]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[18]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[2]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[18]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[2]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[18]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[2])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed2)
);

IOBUF IOBUF_2(
	.I(videosoc_ddrphy_dq_o2),
	.T(videosoc_ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(videosoc_ddrphy_dq_i_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[3]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[19]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[3]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[19]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[3]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[19]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[3]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[19]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o3),
	.TQ(videosoc_ddrphy_dq_t3)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed3),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[19]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[3]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[19]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[3]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[19]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[3]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[19]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[3])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed3)
);

IOBUF IOBUF_3(
	.I(videosoc_ddrphy_dq_o3),
	.T(videosoc_ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(videosoc_ddrphy_dq_i_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[4]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[20]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[4]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[20]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[4]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[20]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[4]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[20]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o4),
	.TQ(videosoc_ddrphy_dq_t4)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed4),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[20]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[4]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[20]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[4]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[20]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[4]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[20]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[4])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed4)
);

IOBUF IOBUF_4(
	.I(videosoc_ddrphy_dq_o4),
	.T(videosoc_ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(videosoc_ddrphy_dq_i_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[5]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[21]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[5]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[21]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[5]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[21]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[5]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[21]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o5),
	.TQ(videosoc_ddrphy_dq_t5)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed5),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[21]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[5]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[21]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[5]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[21]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[5]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[21]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[5])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed5)
);

IOBUF IOBUF_5(
	.I(videosoc_ddrphy_dq_o5),
	.T(videosoc_ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(videosoc_ddrphy_dq_i_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[6]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[22]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[6]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[22]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[6]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[22]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[6]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[22]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o6),
	.TQ(videosoc_ddrphy_dq_t6)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed6),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[22]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[6]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[22]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[6]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[22]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[6]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[22]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[6])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed6)
);

IOBUF IOBUF_6(
	.I(videosoc_ddrphy_dq_o6),
	.T(videosoc_ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(videosoc_ddrphy_dq_i_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[7]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[23]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[7]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[23]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[7]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[23]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[7]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[23]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o7),
	.TQ(videosoc_ddrphy_dq_t7)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed7),
	.RST((sys_rst | (videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[23]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[7]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[23]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[7]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[23]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[7]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[23]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[7])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[0] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed7)
);

IOBUF IOBUF_7(
	.I(videosoc_ddrphy_dq_o7),
	.T(videosoc_ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(videosoc_ddrphy_dq_i_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[8]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[24]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[8]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[24]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[8]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[24]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[8]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[24]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o8),
	.TQ(videosoc_ddrphy_dq_t8)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed8),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[24]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[8]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[24]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[8]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[24]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[8]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[24]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[8])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed8)
);

IOBUF IOBUF_8(
	.I(videosoc_ddrphy_dq_o8),
	.T(videosoc_ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(videosoc_ddrphy_dq_i_nodelay8)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[9]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[25]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[9]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[25]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[9]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[25]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[9]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[25]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o9),
	.TQ(videosoc_ddrphy_dq_t9)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed9),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[25]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[9]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[25]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[9]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[25]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[9]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[25]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[9])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed9)
);

IOBUF IOBUF_9(
	.I(videosoc_ddrphy_dq_o9),
	.T(videosoc_ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(videosoc_ddrphy_dq_i_nodelay9)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[10]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[26]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[10]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[26]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[10]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[26]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[10]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[26]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o10),
	.TQ(videosoc_ddrphy_dq_t10)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed10),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[26]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[10]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[26]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[10]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[26]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[10]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[26]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[10])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed10)
);

IOBUF IOBUF_10(
	.I(videosoc_ddrphy_dq_o10),
	.T(videosoc_ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(videosoc_ddrphy_dq_i_nodelay10)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[11]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[27]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[11]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[27]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[11]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[27]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[11]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[27]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o11),
	.TQ(videosoc_ddrphy_dq_t11)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed11),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[27]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[11]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[27]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[11]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[27]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[11]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[27]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[11])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed11)
);

IOBUF IOBUF_11(
	.I(videosoc_ddrphy_dq_o11),
	.T(videosoc_ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(videosoc_ddrphy_dq_i_nodelay11)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[12]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[28]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[12]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[28]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[12]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[28]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[12]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[28]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o12),
	.TQ(videosoc_ddrphy_dq_t12)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed12),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[28]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[12]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[28]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[12]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[28]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[12]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[28]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[12])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed12)
);

IOBUF IOBUF_12(
	.I(videosoc_ddrphy_dq_o12),
	.T(videosoc_ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(videosoc_ddrphy_dq_i_nodelay12)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[13]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[29]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[13]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[29]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[13]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[29]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[13]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[29]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o13),
	.TQ(videosoc_ddrphy_dq_t13)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed13),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[29]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[13]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[29]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[13]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[29]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[13]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[29]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[13])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed13)
);

IOBUF IOBUF_13(
	.I(videosoc_ddrphy_dq_o13),
	.T(videosoc_ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(videosoc_ddrphy_dq_i_nodelay13)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[14]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[30]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[14]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[30]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[14]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[30]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[14]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[30]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o14),
	.TQ(videosoc_ddrphy_dq_t14)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed14),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[30]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[14]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[30]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[14]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[30]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[14]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[30]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[14])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed14)
);

IOBUF IOBUF_14(
	.I(videosoc_ddrphy_dq_o14),
	.T(videosoc_ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(videosoc_ddrphy_dq_i_nodelay14)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(videosoc_ddrphy_dfi_p0_wrdata[15]),
	.D2(videosoc_ddrphy_dfi_p0_wrdata[31]),
	.D3(videosoc_ddrphy_dfi_p1_wrdata[15]),
	.D4(videosoc_ddrphy_dfi_p1_wrdata[31]),
	.D5(videosoc_ddrphy_dfi_p2_wrdata[15]),
	.D6(videosoc_ddrphy_dfi_p2_wrdata[31]),
	.D7(videosoc_ddrphy_dfi_p3_wrdata[15]),
	.D8(videosoc_ddrphy_dfi_p3_wrdata[31]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(videosoc_ddrphy_dq_o15),
	.TQ(videosoc_ddrphy_dq_t15)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(videosoc_ddrphy_dq_i_delayed15),
	.RST((sys_rst | (videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(videosoc_ddrphy_dfi_p3_rddata[31]),
	.Q2(videosoc_ddrphy_dfi_p3_rddata[15]),
	.Q3(videosoc_ddrphy_dfi_p2_rddata[31]),
	.Q4(videosoc_ddrphy_dfi_p2_rddata[15]),
	.Q5(videosoc_ddrphy_dfi_p1_rddata[31]),
	.Q6(videosoc_ddrphy_dfi_p1_rddata[15]),
	.Q7(videosoc_ddrphy_dfi_p0_rddata[31]),
	.Q8(videosoc_ddrphy_dfi_p0_rddata[15])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(videosoc_ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((videosoc_ddrphy_storage[1] & videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(videosoc_ddrphy_dq_i_delayed15)
);

IOBUF IOBUF_15(
	.I(videosoc_ddrphy_dq_o15),
	.T(videosoc_ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(videosoc_ddrphy_dq_i_nodelay15)
);

reg [24:0] storage_2[0:7];
reg [2:0] memadr_3;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine0_wrport_we)
		storage_2[videosoc_sdram_bankmachine0_wrport_adr] <= videosoc_sdram_bankmachine0_wrport_dat_w;
	memadr_3 <= videosoc_sdram_bankmachine0_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine0_wrport_dat_r = storage_2[memadr_3];
assign videosoc_sdram_bankmachine0_rdport_dat_r = storage_2[videosoc_sdram_bankmachine0_rdport_adr];

reg [24:0] storage_3[0:7];
reg [2:0] memadr_4;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine1_wrport_we)
		storage_3[videosoc_sdram_bankmachine1_wrport_adr] <= videosoc_sdram_bankmachine1_wrport_dat_w;
	memadr_4 <= videosoc_sdram_bankmachine1_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine1_wrport_dat_r = storage_3[memadr_4];
assign videosoc_sdram_bankmachine1_rdport_dat_r = storage_3[videosoc_sdram_bankmachine1_rdport_adr];

reg [24:0] storage_4[0:7];
reg [2:0] memadr_5;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine2_wrport_we)
		storage_4[videosoc_sdram_bankmachine2_wrport_adr] <= videosoc_sdram_bankmachine2_wrport_dat_w;
	memadr_5 <= videosoc_sdram_bankmachine2_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine2_wrport_dat_r = storage_4[memadr_5];
assign videosoc_sdram_bankmachine2_rdport_dat_r = storage_4[videosoc_sdram_bankmachine2_rdport_adr];

reg [24:0] storage_5[0:7];
reg [2:0] memadr_6;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine3_wrport_we)
		storage_5[videosoc_sdram_bankmachine3_wrport_adr] <= videosoc_sdram_bankmachine3_wrport_dat_w;
	memadr_6 <= videosoc_sdram_bankmachine3_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine3_wrport_dat_r = storage_5[memadr_6];
assign videosoc_sdram_bankmachine3_rdport_dat_r = storage_5[videosoc_sdram_bankmachine3_rdport_adr];

reg [24:0] storage_6[0:7];
reg [2:0] memadr_7;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine4_wrport_we)
		storage_6[videosoc_sdram_bankmachine4_wrport_adr] <= videosoc_sdram_bankmachine4_wrport_dat_w;
	memadr_7 <= videosoc_sdram_bankmachine4_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine4_wrport_dat_r = storage_6[memadr_7];
assign videosoc_sdram_bankmachine4_rdport_dat_r = storage_6[videosoc_sdram_bankmachine4_rdport_adr];

reg [24:0] storage_7[0:7];
reg [2:0] memadr_8;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine5_wrport_we)
		storage_7[videosoc_sdram_bankmachine5_wrport_adr] <= videosoc_sdram_bankmachine5_wrport_dat_w;
	memadr_8 <= videosoc_sdram_bankmachine5_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine5_wrport_dat_r = storage_7[memadr_8];
assign videosoc_sdram_bankmachine5_rdport_dat_r = storage_7[videosoc_sdram_bankmachine5_rdport_adr];

reg [24:0] storage_8[0:7];
reg [2:0] memadr_9;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine6_wrport_we)
		storage_8[videosoc_sdram_bankmachine6_wrport_adr] <= videosoc_sdram_bankmachine6_wrport_dat_w;
	memadr_9 <= videosoc_sdram_bankmachine6_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine6_wrport_dat_r = storage_8[memadr_9];
assign videosoc_sdram_bankmachine6_rdport_dat_r = storage_8[videosoc_sdram_bankmachine6_rdport_adr];

reg [24:0] storage_9[0:7];
reg [2:0] memadr_10;
always @(posedge sys_clk) begin
	if (videosoc_sdram_bankmachine7_wrport_we)
		storage_9[videosoc_sdram_bankmachine7_wrport_adr] <= videosoc_sdram_bankmachine7_wrport_dat_w;
	memadr_10 <= videosoc_sdram_bankmachine7_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign videosoc_sdram_bankmachine7_wrport_dat_r = storage_9[memadr_10];
assign videosoc_sdram_bankmachine7_rdport_dat_r = storage_9[videosoc_sdram_bankmachine7_rdport_adr];

reg [23:0] tag_mem[0:511];
reg [8:0] memadr_11;
always @(posedge sys_clk) begin
	if (videosoc_tag_port_we)
		tag_mem[videosoc_tag_port_adr] <= videosoc_tag_port_dat_w;
	memadr_11 <= videosoc_tag_port_adr;
end

assign videosoc_tag_port_dat_r = tag_mem[memadr_11];

STARTUPE2 STARTUPE2(
	.CLK(1'd0),
	.GSR(1'd0),
	.GTS(1'd0),
	.KEYCLEARB(1'd0),
	.PACK(1'd0),
	.USRCCLKO(videosoc_clk0),
	.USRCCLKTS(1'd0),
	.USRDONEO(1'd1),
	.USRDONETS(1'd1)
);

IBUF IBUF(
	.I(eth_clocks_rx),
	.O(ethphy_eth_rx_clk_ibuf)
);

BUFG BUFG_5(
	.I(ethphy_eth_rx_clk_ibuf),
	.O(eth_rx_clk)
);

PLLE2_BASE #(
	.CLKFBOUT_MULT(4'd8),
	.CLKIN1_PERIOD(8.0),
	.CLKOUT0_DIVIDE(4'd8),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(4'd8),
	.CLKOUT1_PHASE(90.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_BASE_1 (
	.CLKFBIN(ethphy_pll_fb),
	.CLKIN1(eth_rx_clk),
	.CLKFBOUT(ethphy_pll_fb),
	.CLKOUT0(ethphy_pll_clk_tx),
	.CLKOUT1(ethphy_pll_clk_tx90),
	.LOCKED(ethphy_pll_locked)
);

BUFG BUFG_6(
	.I(ethphy_pll_clk_tx),
	.O(eth_tx_clk)
);

BUFG BUFG_7(
	.I(ethphy_pll_clk_tx90),
	.O(eth_tx90_clk)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR (
	.C(eth_tx90_clk),
	.CE(1'd1),
	.D1(1'd1),
	.D2(1'd0),
	.R(1'd0),
	.S(1'd0),
	.Q(ethphy_eth_tx_clk_obuf)
);

OBUF OBUF(
	.I(ethphy_eth_tx_clk_obuf),
	.O(eth_clocks_tx)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_1 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(ethphy_sink_valid),
	.D2(ethphy_sink_valid),
	.R(1'd0),
	.S(1'd0),
	.Q(ethphy_tx_ctl_obuf)
);

OBUF OBUF_1(
	.I(ethphy_tx_ctl_obuf),
	.O(eth_tx_ctl)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_2 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(ethphy_sink_payload_data[0]),
	.D2(ethphy_sink_payload_data[4]),
	.R(1'd0),
	.S(1'd0),
	.Q(ethphy_tx_data_obuf[0])
);

OBUF OBUF_2(
	.I(ethphy_tx_data_obuf[0]),
	.O(eth_tx_data[0])
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_3 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(ethphy_sink_payload_data[1]),
	.D2(ethphy_sink_payload_data[5]),
	.R(1'd0),
	.S(1'd0),
	.Q(ethphy_tx_data_obuf[1])
);

OBUF OBUF_3(
	.I(ethphy_tx_data_obuf[1]),
	.O(eth_tx_data[1])
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_4 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(ethphy_sink_payload_data[2]),
	.D2(ethphy_sink_payload_data[6]),
	.R(1'd0),
	.S(1'd0),
	.Q(ethphy_tx_data_obuf[2])
);

OBUF OBUF_4(
	.I(ethphy_tx_data_obuf[2]),
	.O(eth_tx_data[2])
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_5 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(ethphy_sink_payload_data[3]),
	.D2(ethphy_sink_payload_data[7]),
	.R(1'd0),
	.S(1'd0),
	.Q(ethphy_tx_data_obuf[3])
);

OBUF OBUF_5(
	.I(ethphy_tx_data_obuf[3]),
	.O(eth_tx_data[3])
);

IBUF IBUF_1(
	.I(eth_rx_ctl),
	.O(ethphy_rx_ctl_ibuf)
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_16 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(ethphy_rx_ctl_ibuf),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(ethphy_rx_ctl_idelay)
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(ethphy_rx_ctl_idelay),
	.R(1'd0),
	.S(1'd0),
	.Q1(ethphy_rx_ctl)
);

IBUF IBUF_2(
	.I(eth_rx_data[0]),
	.O(ethphy_rx_data_ibuf[0])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_17 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(ethphy_rx_data_ibuf[0]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(ethphy_rx_data_idelay[0])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_1 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(ethphy_rx_data_idelay[0]),
	.R(1'd0),
	.S(1'd0),
	.Q1(ethphy_rx_data[0]),
	.Q2(ethphy_rx_data[4])
);

IBUF IBUF_3(
	.I(eth_rx_data[1]),
	.O(ethphy_rx_data_ibuf[1])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_18 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(ethphy_rx_data_ibuf[1]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(ethphy_rx_data_idelay[1])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_2 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(ethphy_rx_data_idelay[1]),
	.R(1'd0),
	.S(1'd0),
	.Q1(ethphy_rx_data[1]),
	.Q2(ethphy_rx_data[5])
);

IBUF IBUF_4(
	.I(eth_rx_data[2]),
	.O(ethphy_rx_data_ibuf[2])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_19 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(ethphy_rx_data_ibuf[2]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(ethphy_rx_data_idelay[2])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_3 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(ethphy_rx_data_idelay[2]),
	.R(1'd0),
	.S(1'd0),
	.Q1(ethphy_rx_data[2]),
	.Q2(ethphy_rx_data[6])
);

IBUF IBUF_5(
	.I(eth_rx_data[3]),
	.O(ethphy_rx_data_ibuf[3])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_20 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(ethphy_rx_data_ibuf[3]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(ethphy_rx_data_idelay[3])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_4 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(ethphy_rx_data_idelay[3]),
	.R(1'd0),
	.S(1'd0),
	.Q1(ethphy_rx_data[3]),
	.Q2(ethphy_rx_data[7])
);

assign eth_mdio = ethphy_data_oe ? ethphy_data_w : 1'bz;
assign ethphy_data_r = eth_mdio;

reg [11:0] storage_10[0:4];
reg [2:0] memadr_12;
always @(posedge eth_rx_clk) begin
	if (ethmac_crc32_checker_syncfifo_wrport_we)
		storage_10[ethmac_crc32_checker_syncfifo_wrport_adr] <= ethmac_crc32_checker_syncfifo_wrport_dat_w;
	memadr_12 <= ethmac_crc32_checker_syncfifo_wrport_adr;
end

always @(posedge eth_rx_clk) begin
end

assign ethmac_crc32_checker_syncfifo_wrport_dat_r = storage_10[memadr_12];
assign ethmac_crc32_checker_syncfifo_rdport_dat_r = storage_10[ethmac_crc32_checker_syncfifo_rdport_adr];

reg [41:0] storage_11[0:63];
reg [5:0] memadr_13;
reg [41:0] memdat_2;
always @(posedge sys_clk) begin
	if (ethmac_tx_cdc_wrport_we)
		storage_11[ethmac_tx_cdc_wrport_adr] <= ethmac_tx_cdc_wrport_dat_w;
	memadr_13 <= ethmac_tx_cdc_wrport_adr;
end

always @(posedge eth_tx_clk) begin
	memdat_2 <= storage_11[ethmac_tx_cdc_rdport_adr];
end

assign ethmac_tx_cdc_wrport_dat_r = storage_11[memadr_13];
assign ethmac_tx_cdc_rdport_dat_r = memdat_2;

reg [41:0] storage_12[0:63];
reg [5:0] memadr_14;
reg [41:0] memdat_3;
always @(posedge eth_rx_clk) begin
	if (ethmac_rx_cdc_wrport_we)
		storage_12[ethmac_rx_cdc_wrport_adr] <= ethmac_rx_cdc_wrport_dat_w;
	memadr_14 <= ethmac_rx_cdc_wrport_adr;
end

always @(posedge sys_clk) begin
	memdat_3 <= storage_12[ethmac_rx_cdc_rdport_adr];
end

assign ethmac_rx_cdc_wrport_dat_r = storage_12[memadr_14];
assign ethmac_rx_cdc_rdport_dat_r = memdat_3;

reg [34:0] storage_13[0:1];
reg [0:0] memadr_15;
always @(posedge sys_clk) begin
	if (ethmac_writer_fifo_wrport_we)
		storage_13[ethmac_writer_fifo_wrport_adr] <= ethmac_writer_fifo_wrport_dat_w;
	memadr_15 <= ethmac_writer_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign ethmac_writer_fifo_wrport_dat_r = storage_13[memadr_15];
assign ethmac_writer_fifo_rdport_dat_r = storage_13[ethmac_writer_fifo_rdport_adr];

reg [31:0] mem_3[0:381];
reg [8:0] memadr_16;
reg [31:0] memdat_4;
always @(posedge sys_clk) begin
	if (ethmac_writer_memory0_we)
		mem_3[ethmac_writer_memory0_adr] <= ethmac_writer_memory0_dat_w;
	memadr_16 <= ethmac_writer_memory0_adr;
end

always @(posedge sys_clk) begin
	memdat_4 <= mem_3[ethmac_sram0_adr0];
end

assign ethmac_writer_memory0_dat_r = mem_3[memadr_16];
assign ethmac_sram0_dat_r0 = memdat_4;

reg [31:0] mem_4[0:381];
reg [8:0] memadr_17;
reg [31:0] memdat_5;
always @(posedge sys_clk) begin
	if (ethmac_writer_memory1_we)
		mem_4[ethmac_writer_memory1_adr] <= ethmac_writer_memory1_dat_w;
	memadr_17 <= ethmac_writer_memory1_adr;
end

always @(posedge sys_clk) begin
	memdat_5 <= mem_4[ethmac_sram1_adr0];
end

assign ethmac_writer_memory1_dat_r = mem_4[memadr_17];
assign ethmac_sram1_dat_r0 = memdat_5;

reg [13:0] storage_14[0:1];
reg [0:0] memadr_18;
always @(posedge sys_clk) begin
	if (ethmac_reader_fifo_wrport_we)
		storage_14[ethmac_reader_fifo_wrport_adr] <= ethmac_reader_fifo_wrport_dat_w;
	memadr_18 <= ethmac_reader_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign ethmac_reader_fifo_wrport_dat_r = storage_14[memadr_18];
assign ethmac_reader_fifo_rdport_dat_r = storage_14[ethmac_reader_fifo_rdport_adr];

reg [7:0] edid_mem[0:127];
reg [7:0] memdat_6;
reg [6:0] memadr_19;
always @(posedge sys_clk) begin
	memdat_6 <= edid_mem[edid_adr];
end

always @(posedge sys_clk) begin
	if (videosoc_sram0_we)
		edid_mem[videosoc_sram0_adr] <= videosoc_sram0_dat_w;
	memadr_19 <= videosoc_sram0_adr;
end

assign edid_dat_r = memdat_6;
assign videosoc_sram0_dat_r = edid_mem[memadr_19];

initial begin
	$readmemh("edid_mem.init", edid_mem);
end

assign hdmi_in_sda = edid_sda_drv_reg ? 1'd0 : 1'bz;
assign edid_sda_i_async = hdmi_in_sda;

IBUFDS hdmi_in_ibufds(
	.I(hdmi_in_clk_p),
	.IB(hdmi_in_clk_n),
	.O(clk_input)
);

BUFG BUFG_8(
	.I(clk_input),
	.O(clk_input_bufg)
);

MMCME2_ADV #(
	.BANDWIDTH("OPTIMIZED"),
	.CLKFBOUT_MULT_F(10.0),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(6.734006734006734),
	.CLKOUT0_DIVIDE_F(4'd10),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(4'd8),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(2'd2),
	.CLKOUT2_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01)
) MMCME2_ADV (
	.CLKFBIN(mmcm_fb),
	.CLKIN1(clk_input),
	.DADDR(mmcm_adr_storage),
	.DCLK(sys_clk),
	.DEN((mmcm_read_re | mmcm_write_re)),
	.DI(mmcm_dat_w_storage),
	.DWE(mmcm_write_re),
	.RST(mmcm_reset_storage),
	.CLKFBOUT(mmcm_fb),
	.CLKOUT0(mmcm_clk0),
	.CLKOUT1(mmcm_clk1),
	.CLKOUT2(mmcm_clk2),
	.DO(mmcm_dat_r_status),
	.DRDY(mmcm_drdy),
	.LOCKED(mmcm_locked)
);

BUFG BUFG_9(
	.I(mmcm_clk0),
	.O(hdmi_in0_pix_clk)
);

BUFR BUFR(
	.I(mmcm_clk1),
	.O(pix1p25x_clk)
);

BUFIO BUFIO(
	.I(mmcm_clk2),
	.O(hdmi_in0_pix5x_clk)
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT(
	.I(hdmi_in_data0_p),
	.IB(hdmi_in_data0_n),
	.O(s7datacapture0_serdes_m_i_nodelay),
	.OB(s7datacapture0_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_21 (
	.C(pix1p25x_clk),
	.CE(s7datacapture0_delay_master_ce),
	.IDATAIN(s7datacapture0_serdes_m_i_nodelay),
	.INC(s7datacapture0_delay_master_inc),
	.LD(s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(s7datacapture0_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_16 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(s7datacapture0_serdes_m_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(s7datacapture0_serdes_m_q[7]),
	.Q2(s7datacapture0_serdes_m_q[6]),
	.Q3(s7datacapture0_serdes_m_q[5]),
	.Q4(s7datacapture0_serdes_m_q[4]),
	.Q5(s7datacapture0_serdes_m_q[3]),
	.Q6(s7datacapture0_serdes_m_q[2]),
	.Q7(s7datacapture0_serdes_m_q[1]),
	.Q8(s7datacapture0_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_22 (
	.C(pix1p25x_clk),
	.CE(s7datacapture0_delay_slave_ce),
	.IDATAIN(s7datacapture0_serdes_s_i_nodelay),
	.INC(s7datacapture0_delay_slave_inc),
	.LD(s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(s7datacapture0_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_17 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(s7datacapture0_serdes_s_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(s7datacapture0_serdes_s_q[7]),
	.Q2(s7datacapture0_serdes_s_q[6]),
	.Q3(s7datacapture0_serdes_s_q[5]),
	.Q4(s7datacapture0_serdes_s_q[4]),
	.Q5(s7datacapture0_serdes_s_q[3]),
	.Q6(s7datacapture0_serdes_s_q[2]),
	.Q7(s7datacapture0_serdes_s_q[1]),
	.Q8(s7datacapture0_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_1(
	.I(hdmi_in_data1_p),
	.IB(hdmi_in_data1_n),
	.O(s7datacapture1_serdes_m_i_nodelay),
	.OB(s7datacapture1_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_23 (
	.C(pix1p25x_clk),
	.CE(s7datacapture1_delay_master_ce),
	.IDATAIN(s7datacapture1_serdes_m_i_nodelay),
	.INC(s7datacapture1_delay_master_inc),
	.LD(s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(s7datacapture1_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_18 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(s7datacapture1_serdes_m_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(s7datacapture1_serdes_m_q[7]),
	.Q2(s7datacapture1_serdes_m_q[6]),
	.Q3(s7datacapture1_serdes_m_q[5]),
	.Q4(s7datacapture1_serdes_m_q[4]),
	.Q5(s7datacapture1_serdes_m_q[3]),
	.Q6(s7datacapture1_serdes_m_q[2]),
	.Q7(s7datacapture1_serdes_m_q[1]),
	.Q8(s7datacapture1_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_24 (
	.C(pix1p25x_clk),
	.CE(s7datacapture1_delay_slave_ce),
	.IDATAIN(s7datacapture1_serdes_s_i_nodelay),
	.INC(s7datacapture1_delay_slave_inc),
	.LD(s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(s7datacapture1_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_19 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(s7datacapture1_serdes_s_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(s7datacapture1_serdes_s_q[7]),
	.Q2(s7datacapture1_serdes_s_q[6]),
	.Q3(s7datacapture1_serdes_s_q[5]),
	.Q4(s7datacapture1_serdes_s_q[4]),
	.Q5(s7datacapture1_serdes_s_q[3]),
	.Q6(s7datacapture1_serdes_s_q[2]),
	.Q7(s7datacapture1_serdes_s_q[1]),
	.Q8(s7datacapture1_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_2(
	.I(hdmi_in_data2_p),
	.IB(hdmi_in_data2_n),
	.O(s7datacapture2_serdes_m_i_nodelay),
	.OB(s7datacapture2_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_25 (
	.C(pix1p25x_clk),
	.CE(s7datacapture2_delay_master_ce),
	.IDATAIN(s7datacapture2_serdes_m_i_nodelay),
	.INC(s7datacapture2_delay_master_inc),
	.LD(s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(s7datacapture2_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_20 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(s7datacapture2_serdes_m_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(s7datacapture2_serdes_m_q[7]),
	.Q2(s7datacapture2_serdes_m_q[6]),
	.Q3(s7datacapture2_serdes_m_q[5]),
	.Q4(s7datacapture2_serdes_m_q[4]),
	.Q5(s7datacapture2_serdes_m_q[3]),
	.Q6(s7datacapture2_serdes_m_q[2]),
	.Q7(s7datacapture2_serdes_m_q[1]),
	.Q8(s7datacapture2_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_26 (
	.C(pix1p25x_clk),
	.CE(s7datacapture2_delay_slave_ce),
	.IDATAIN(s7datacapture2_serdes_s_i_nodelay),
	.INC(s7datacapture2_delay_slave_inc),
	.LD(s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(s7datacapture2_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_21 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(s7datacapture2_serdes_s_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(s7datacapture2_serdes_s_q[7]),
	.Q2(s7datacapture2_serdes_s_q[6]),
	.Q3(s7datacapture2_serdes_s_q[5]),
	.Q4(s7datacapture2_serdes_s_q[4]),
	.Q5(s7datacapture2_serdes_s_q[3]),
	.Q6(s7datacapture2_serdes_s_q[2]),
	.Q7(s7datacapture2_serdes_s_q[1]),
	.Q8(s7datacapture2_serdes_s_q[0])
);

reg [10:0] storage_15[0:7];
reg [2:0] memadr_20;
always @(posedge hdmi_in0_pix_clk) begin
	if (chansync_syncbuffer0_wrport_we)
		storage_15[chansync_syncbuffer0_wrport_adr] <= chansync_syncbuffer0_wrport_dat_w;
	memadr_20 <= chansync_syncbuffer0_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign chansync_syncbuffer0_wrport_dat_r = storage_15[memadr_20];
assign chansync_syncbuffer0_rdport_dat_r = storage_15[chansync_syncbuffer0_rdport_adr];

reg [10:0] storage_16[0:7];
reg [2:0] memadr_21;
always @(posedge hdmi_in0_pix_clk) begin
	if (chansync_syncbuffer1_wrport_we)
		storage_16[chansync_syncbuffer1_wrport_adr] <= chansync_syncbuffer1_wrport_dat_w;
	memadr_21 <= chansync_syncbuffer1_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign chansync_syncbuffer1_wrport_dat_r = storage_16[memadr_21];
assign chansync_syncbuffer1_rdport_dat_r = storage_16[chansync_syncbuffer1_rdport_adr];

reg [10:0] storage_17[0:7];
reg [2:0] memadr_22;
always @(posedge hdmi_in0_pix_clk) begin
	if (chansync_syncbuffer2_wrport_we)
		storage_17[chansync_syncbuffer2_wrport_adr] <= chansync_syncbuffer2_wrport_dat_w;
	memadr_22 <= chansync_syncbuffer2_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign chansync_syncbuffer2_wrport_dat_r = storage_17[memadr_22];
assign chansync_syncbuffer2_rdport_dat_r = storage_17[chansync_syncbuffer2_rdport_adr];

reg [130:0] storage_18[0:511];
reg [8:0] memadr_23;
reg [130:0] memdat_7;
always @(posedge hdmi_in0_pix_clk) begin
	if (frame_fifo_wrport_we)
		storage_18[frame_fifo_wrport_adr] <= frame_fifo_wrport_dat_w;
	memadr_23 <= frame_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memdat_7 <= storage_18[frame_fifo_rdport_adr];
end

assign frame_fifo_wrport_dat_r = storage_18[memadr_23];
assign frame_fifo_rdport_dat_r = memdat_7;

reg [129:0] storage_19[0:15];
reg [3:0] memadr_24;
always @(posedge sys_clk) begin
	if (dma_fifo_wrport_we)
		storage_19[dma_fifo_wrport_adr] <= dma_fifo_wrport_dat_w;
	memadr_24 <= dma_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign dma_fifo_wrport_dat_r = storage_19[memadr_24];
assign dma_fifo_rdport_dat_r = storage_19[dma_fifo_rdport_adr];

reg [27:0] storage_20[0:3];
reg [1:0] memadr_25;
reg [27:0] memdat_8;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi_out0_dram_port_cmd_fifo_wrport_we)
		storage_20[hdmi_out0_dram_port_cmd_fifo_wrport_adr] <= hdmi_out0_dram_port_cmd_fifo_wrport_dat_w;
	memadr_25 <= hdmi_out0_dram_port_cmd_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memdat_8 <= storage_20[hdmi_out0_dram_port_cmd_fifo_rdport_adr];
end

assign hdmi_out0_dram_port_cmd_fifo_wrport_dat_r = storage_20[memadr_25];
assign hdmi_out0_dram_port_cmd_fifo_rdport_dat_r = memdat_8;

reg [129:0] storage_21[0:15];
reg [3:0] memadr_26;
reg [129:0] memdat_9;
always @(posedge sys_clk) begin
	if (hdmi_out0_dram_port_rdata_fifo_wrport_we)
		storage_21[hdmi_out0_dram_port_rdata_fifo_wrport_adr] <= hdmi_out0_dram_port_rdata_fifo_wrport_dat_w;
	memadr_26 <= hdmi_out0_dram_port_rdata_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	memdat_9 <= storage_21[hdmi_out0_dram_port_rdata_fifo_rdport_adr];
end

assign hdmi_out0_dram_port_rdata_fifo_wrport_dat_r = storage_21[memadr_26];
assign hdmi_out0_dram_port_rdata_fifo_rdport_dat_r = memdat_9;

reg [9:0] storage_22[0:3];
reg [1:0] memadr_27;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi_out0_dram_port_cmd_buffer_wrport_we)
		storage_22[hdmi_out0_dram_port_cmd_buffer_wrport_adr] <= hdmi_out0_dram_port_cmd_buffer_wrport_dat_w;
	memadr_27 <= hdmi_out0_dram_port_cmd_buffer_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi_out0_dram_port_cmd_buffer_wrport_dat_r = storage_22[memadr_27];
assign hdmi_out0_dram_port_cmd_buffer_rdport_dat_r = storage_22[hdmi_out0_dram_port_cmd_buffer_rdport_adr];

reg [161:0] storage_23[0:1];
reg [0:0] memadr_28;
reg [161:0] memdat_10;
always @(posedge sys_clk) begin
	if (hdmi_out0_core_initiator_cdc_wrport_we)
		storage_23[hdmi_out0_core_initiator_cdc_wrport_adr] <= hdmi_out0_core_initiator_cdc_wrport_dat_w;
	memadr_28 <= hdmi_out0_core_initiator_cdc_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	memdat_10 <= storage_23[hdmi_out0_core_initiator_cdc_rdport_adr];
end

assign hdmi_out0_core_initiator_cdc_wrport_dat_r = storage_23[memadr_28];
assign hdmi_out0_core_initiator_cdc_rdport_dat_r = memdat_10;

reg [17:0] storage_24[0:4095];
reg [11:0] memadr_29;
reg [17:0] memdat_11;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi_out0_core_dmareader_fifo_wrport_we)
		storage_24[hdmi_out0_core_dmareader_fifo_wrport_adr] <= hdmi_out0_core_dmareader_fifo_wrport_dat_w;
	memadr_29 <= hdmi_out0_core_dmareader_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi_out0_core_dmareader_fifo_rdport_re)
		memdat_11 <= storage_24[hdmi_out0_core_dmareader_fifo_rdport_adr];
end

assign hdmi_out0_core_dmareader_fifo_wrport_dat_r = storage_24[memadr_29];
assign hdmi_out0_core_dmareader_fifo_rdport_dat_r = memdat_11;

MMCME2_ADV #(
	.BANDWIDTH("OPTIMIZED"),
	.CLKFBOUT_MULT_F(30.0),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(10.0),
	.CLKOUT0_DIVIDE_F(10.0),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(2'd2),
	.CLKOUT1_PHASE(0.0),
	.DIVCLK_DIVIDE(2'd2),
	.REF_JITTER1(0.01)
) MMCME2_ADV_1 (
	.CLKFBIN(hdmi_out0_driver_s7hdmioutclocking_mmcm_fb),
	.CLKIN1(clk100_clk),
	.DADDR(hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage),
	.DCLK(sys_clk),
	.DEN((hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re | hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re)),
	.DI(hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage),
	.DWE(hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re),
	.RST(hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage),
	.CLKFBOUT(hdmi_out0_driver_s7hdmioutclocking_mmcm_fb),
	.CLKOUT0(hdmi_out0_driver_s7hdmioutclocking_mmcm_clk0),
	.CLKOUT1(hdmi_out0_driver_s7hdmioutclocking_mmcm_clk1),
	.DO(hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status),
	.DRDY(hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy),
	.LOCKED(hdmi_out0_driver_s7hdmioutclocking_mmcm_locked)
);

BUFG BUFG_10(
	.I(hdmi_out0_driver_s7hdmioutclocking_mmcm_clk0),
	.O(hdmi_out0_pix_clk)
);

BUFG BUFG_11(
	.I(hdmi_out0_driver_s7hdmioutclocking_mmcm_clk1),
	.O(hdmi_out0_pix5x_clk)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_45 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(hdmi_out0_driver_s7hdmioutclocking_data1[0]),
	.D2(hdmi_out0_driver_s7hdmioutclocking_data1[1]),
	.D3(hdmi_out0_driver_s7hdmioutclocking_data1[2]),
	.D4(hdmi_out0_driver_s7hdmioutclocking_data1[3]),
	.D5(hdmi_out0_driver_s7hdmioutclocking_data1[4]),
	.D6(hdmi_out0_driver_s7hdmioutclocking_data1[5]),
	.D7(hdmi_out0_driver_s7hdmioutclocking_data1[6]),
	.D8(hdmi_out0_driver_s7hdmioutclocking_data1[7]),
	.OCE(hdmi_out0_driver_s7hdmioutclocking_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(hdmi_out0_driver_s7hdmioutclocking_shift[0]),
	.SHIFTIN2(hdmi_out0_driver_s7hdmioutclocking_shift[1]),
	.TCE(1'd0),
	.OQ(hdmi_out0_driver_s7hdmioutclocking_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_46 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(hdmi_out0_driver_s7hdmioutclocking_data1[8]),
	.D4(hdmi_out0_driver_s7hdmioutclocking_data1[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(hdmi_out0_driver_s7hdmioutclocking_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(hdmi_out0_driver_s7hdmioutclocking_shift[0]),
	.SHIFTOUT2(hdmi_out0_driver_s7hdmioutclocking_shift[1])
);

OBUFDS OBUFDS_1(
	.I(hdmi_out0_driver_s7hdmioutclocking_pad_se),
	.O(hdmi_out_clk_p),
	.OB(hdmi_out_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_47 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(hdmi_out0_driver_hdmi_phy_es0_data[0]),
	.D2(hdmi_out0_driver_hdmi_phy_es0_data[1]),
	.D3(hdmi_out0_driver_hdmi_phy_es0_data[2]),
	.D4(hdmi_out0_driver_hdmi_phy_es0_data[3]),
	.D5(hdmi_out0_driver_hdmi_phy_es0_data[4]),
	.D6(hdmi_out0_driver_hdmi_phy_es0_data[5]),
	.D7(hdmi_out0_driver_hdmi_phy_es0_data[6]),
	.D8(hdmi_out0_driver_hdmi_phy_es0_data[7]),
	.OCE(hdmi_out0_driver_hdmi_phy_es0_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(hdmi_out0_driver_hdmi_phy_es0_shift[0]),
	.SHIFTIN2(hdmi_out0_driver_hdmi_phy_es0_shift[1]),
	.TCE(1'd0),
	.OQ(hdmi_out0_driver_hdmi_phy_es0_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_48 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(hdmi_out0_driver_hdmi_phy_es0_data[8]),
	.D4(hdmi_out0_driver_hdmi_phy_es0_data[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(hdmi_out0_driver_hdmi_phy_es0_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(hdmi_out0_driver_hdmi_phy_es0_shift[0]),
	.SHIFTOUT2(hdmi_out0_driver_hdmi_phy_es0_shift[1])
);

OBUFDS OBUFDS_2(
	.I(hdmi_out0_driver_hdmi_phy_es0_pad_se),
	.O(hdmi_out_data0_p),
	.OB(hdmi_out_data0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_49 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(hdmi_out0_driver_hdmi_phy_es1_data[0]),
	.D2(hdmi_out0_driver_hdmi_phy_es1_data[1]),
	.D3(hdmi_out0_driver_hdmi_phy_es1_data[2]),
	.D4(hdmi_out0_driver_hdmi_phy_es1_data[3]),
	.D5(hdmi_out0_driver_hdmi_phy_es1_data[4]),
	.D6(hdmi_out0_driver_hdmi_phy_es1_data[5]),
	.D7(hdmi_out0_driver_hdmi_phy_es1_data[6]),
	.D8(hdmi_out0_driver_hdmi_phy_es1_data[7]),
	.OCE(hdmi_out0_driver_hdmi_phy_es1_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(hdmi_out0_driver_hdmi_phy_es1_shift[0]),
	.SHIFTIN2(hdmi_out0_driver_hdmi_phy_es1_shift[1]),
	.TCE(1'd0),
	.OQ(hdmi_out0_driver_hdmi_phy_es1_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_50 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(hdmi_out0_driver_hdmi_phy_es1_data[8]),
	.D4(hdmi_out0_driver_hdmi_phy_es1_data[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(hdmi_out0_driver_hdmi_phy_es1_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(hdmi_out0_driver_hdmi_phy_es1_shift[0]),
	.SHIFTOUT2(hdmi_out0_driver_hdmi_phy_es1_shift[1])
);

OBUFDS OBUFDS_3(
	.I(hdmi_out0_driver_hdmi_phy_es1_pad_se),
	.O(hdmi_out_data1_p),
	.OB(hdmi_out_data1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_51 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(hdmi_out0_driver_hdmi_phy_es2_data[0]),
	.D2(hdmi_out0_driver_hdmi_phy_es2_data[1]),
	.D3(hdmi_out0_driver_hdmi_phy_es2_data[2]),
	.D4(hdmi_out0_driver_hdmi_phy_es2_data[3]),
	.D5(hdmi_out0_driver_hdmi_phy_es2_data[4]),
	.D6(hdmi_out0_driver_hdmi_phy_es2_data[5]),
	.D7(hdmi_out0_driver_hdmi_phy_es2_data[6]),
	.D8(hdmi_out0_driver_hdmi_phy_es2_data[7]),
	.OCE(hdmi_out0_driver_hdmi_phy_es2_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(hdmi_out0_driver_hdmi_phy_es2_shift[0]),
	.SHIFTIN2(hdmi_out0_driver_hdmi_phy_es2_shift[1]),
	.TCE(1'd0),
	.OQ(hdmi_out0_driver_hdmi_phy_es2_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_52 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(hdmi_out0_driver_hdmi_phy_es2_data[8]),
	.D4(hdmi_out0_driver_hdmi_phy_es2_data[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(hdmi_out0_driver_hdmi_phy_es2_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(hdmi_out0_driver_hdmi_phy_es2_shift[0]),
	.SHIFTOUT2(hdmi_out0_driver_hdmi_phy_es2_shift[1])
);

OBUFDS OBUFDS_4(
	.I(hdmi_out0_driver_hdmi_phy_es2_pad_se),
	.O(hdmi_out_data2_p),
	.OB(hdmi_out_data2_n)
);

reg [9:0] storage_25[0:3];
reg [1:0] memadr_30;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi_out0_resetinserter_y_fifo_wrport_we)
		storage_25[hdmi_out0_resetinserter_y_fifo_wrport_adr] <= hdmi_out0_resetinserter_y_fifo_wrport_dat_w;
	memadr_30 <= hdmi_out0_resetinserter_y_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi_out0_resetinserter_y_fifo_wrport_dat_r = storage_25[memadr_30];
assign hdmi_out0_resetinserter_y_fifo_rdport_dat_r = storage_25[hdmi_out0_resetinserter_y_fifo_rdport_adr];

reg [9:0] storage_26[0:3];
reg [1:0] memadr_31;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi_out0_resetinserter_cb_fifo_wrport_we)
		storage_26[hdmi_out0_resetinserter_cb_fifo_wrport_adr] <= hdmi_out0_resetinserter_cb_fifo_wrport_dat_w;
	memadr_31 <= hdmi_out0_resetinserter_cb_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi_out0_resetinserter_cb_fifo_wrport_dat_r = storage_26[memadr_31];
assign hdmi_out0_resetinserter_cb_fifo_rdport_dat_r = storage_26[hdmi_out0_resetinserter_cb_fifo_rdport_adr];

reg [9:0] storage_27[0:3];
reg [1:0] memadr_32;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi_out0_resetinserter_cr_fifo_wrport_we)
		storage_27[hdmi_out0_resetinserter_cr_fifo_wrport_adr] <= hdmi_out0_resetinserter_cr_fifo_wrport_dat_w;
	memadr_32 <= hdmi_out0_resetinserter_cr_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi_out0_resetinserter_cr_fifo_wrport_dat_r = storage_27[memadr_32];
assign hdmi_out0_resetinserter_cr_fifo_rdport_dat_r = storage_27[hdmi_out0_resetinserter_cr_fifo_rdport_adr];

reg [7:0] data_mem_grain0[0:511];
reg [8:0] memadr_33;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[0])
		data_mem_grain0[videosoc_data_port_adr] <= videosoc_data_port_dat_w[7:0];
	memadr_33 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[7:0] = data_mem_grain0[memadr_33];

reg [7:0] data_mem_grain1[0:511];
reg [8:0] memadr_34;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[1])
		data_mem_grain1[videosoc_data_port_adr] <= videosoc_data_port_dat_w[15:8];
	memadr_34 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[15:8] = data_mem_grain1[memadr_34];

reg [7:0] data_mem_grain2[0:511];
reg [8:0] memadr_35;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[2])
		data_mem_grain2[videosoc_data_port_adr] <= videosoc_data_port_dat_w[23:16];
	memadr_35 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[23:16] = data_mem_grain2[memadr_35];

reg [7:0] data_mem_grain3[0:511];
reg [8:0] memadr_36;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[3])
		data_mem_grain3[videosoc_data_port_adr] <= videosoc_data_port_dat_w[31:24];
	memadr_36 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[31:24] = data_mem_grain3[memadr_36];

reg [7:0] data_mem_grain4[0:511];
reg [8:0] memadr_37;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[4])
		data_mem_grain4[videosoc_data_port_adr] <= videosoc_data_port_dat_w[39:32];
	memadr_37 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[39:32] = data_mem_grain4[memadr_37];

reg [7:0] data_mem_grain5[0:511];
reg [8:0] memadr_38;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[5])
		data_mem_grain5[videosoc_data_port_adr] <= videosoc_data_port_dat_w[47:40];
	memadr_38 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[47:40] = data_mem_grain5[memadr_38];

reg [7:0] data_mem_grain6[0:511];
reg [8:0] memadr_39;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[6])
		data_mem_grain6[videosoc_data_port_adr] <= videosoc_data_port_dat_w[55:48];
	memadr_39 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[55:48] = data_mem_grain6[memadr_39];

reg [7:0] data_mem_grain7[0:511];
reg [8:0] memadr_40;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[7])
		data_mem_grain7[videosoc_data_port_adr] <= videosoc_data_port_dat_w[63:56];
	memadr_40 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[63:56] = data_mem_grain7[memadr_40];

reg [7:0] data_mem_grain8[0:511];
reg [8:0] memadr_41;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[8])
		data_mem_grain8[videosoc_data_port_adr] <= videosoc_data_port_dat_w[71:64];
	memadr_41 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[71:64] = data_mem_grain8[memadr_41];

reg [7:0] data_mem_grain9[0:511];
reg [8:0] memadr_42;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[9])
		data_mem_grain9[videosoc_data_port_adr] <= videosoc_data_port_dat_w[79:72];
	memadr_42 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[79:72] = data_mem_grain9[memadr_42];

reg [7:0] data_mem_grain10[0:511];
reg [8:0] memadr_43;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[10])
		data_mem_grain10[videosoc_data_port_adr] <= videosoc_data_port_dat_w[87:80];
	memadr_43 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[87:80] = data_mem_grain10[memadr_43];

reg [7:0] data_mem_grain11[0:511];
reg [8:0] memadr_44;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[11])
		data_mem_grain11[videosoc_data_port_adr] <= videosoc_data_port_dat_w[95:88];
	memadr_44 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[95:88] = data_mem_grain11[memadr_44];

reg [7:0] data_mem_grain12[0:511];
reg [8:0] memadr_45;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[12])
		data_mem_grain12[videosoc_data_port_adr] <= videosoc_data_port_dat_w[103:96];
	memadr_45 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[103:96] = data_mem_grain12[memadr_45];

reg [7:0] data_mem_grain13[0:511];
reg [8:0] memadr_46;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[13])
		data_mem_grain13[videosoc_data_port_adr] <= videosoc_data_port_dat_w[111:104];
	memadr_46 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[111:104] = data_mem_grain13[memadr_46];

reg [7:0] data_mem_grain14[0:511];
reg [8:0] memadr_47;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[14])
		data_mem_grain14[videosoc_data_port_adr] <= videosoc_data_port_dat_w[119:112];
	memadr_47 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[119:112] = data_mem_grain14[memadr_47];

reg [7:0] data_mem_grain15[0:511];
reg [8:0] memadr_48;
always @(posedge sys_clk) begin
	if (videosoc_data_port_we[15])
		data_mem_grain15[videosoc_data_port_adr] <= videosoc_data_port_dat_w[127:120];
	memadr_48 <= videosoc_data_port_adr;
end

assign videosoc_data_port_dat_r[127:120] = data_mem_grain15[memadr_48];

reg [7:0] mem_grain0[0:381];
reg [7:0] memdat_12;
reg [8:0] memadr_49;
always @(posedge sys_clk) begin
	memdat_12 <= mem_grain0[ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram0_we[0])
		mem_grain0[ethmac_sram0_adr1] <= ethmac_sram0_dat_w[7:0];
	memadr_49 <= ethmac_sram0_adr1;
end

assign ethmac_reader_memory0_dat_r[7:0] = memdat_12;
assign ethmac_sram0_dat_r1[7:0] = mem_grain0[memadr_49];

reg [7:0] mem_grain1[0:381];
reg [7:0] memdat_13;
reg [8:0] memadr_50;
always @(posedge sys_clk) begin
	memdat_13 <= mem_grain1[ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram0_we[1])
		mem_grain1[ethmac_sram0_adr1] <= ethmac_sram0_dat_w[15:8];
	memadr_50 <= ethmac_sram0_adr1;
end

assign ethmac_reader_memory0_dat_r[15:8] = memdat_13;
assign ethmac_sram0_dat_r1[15:8] = mem_grain1[memadr_50];

reg [7:0] mem_grain2[0:381];
reg [7:0] memdat_14;
reg [8:0] memadr_51;
always @(posedge sys_clk) begin
	memdat_14 <= mem_grain2[ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram0_we[2])
		mem_grain2[ethmac_sram0_adr1] <= ethmac_sram0_dat_w[23:16];
	memadr_51 <= ethmac_sram0_adr1;
end

assign ethmac_reader_memory0_dat_r[23:16] = memdat_14;
assign ethmac_sram0_dat_r1[23:16] = mem_grain2[memadr_51];

reg [7:0] mem_grain3[0:381];
reg [7:0] memdat_15;
reg [8:0] memadr_52;
always @(posedge sys_clk) begin
	memdat_15 <= mem_grain3[ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram0_we[3])
		mem_grain3[ethmac_sram0_adr1] <= ethmac_sram0_dat_w[31:24];
	memadr_52 <= ethmac_sram0_adr1;
end

assign ethmac_reader_memory0_dat_r[31:24] = memdat_15;
assign ethmac_sram0_dat_r1[31:24] = mem_grain3[memadr_52];

reg [7:0] mem_grain0_1[0:381];
reg [7:0] memdat_16;
reg [8:0] memadr_53;
always @(posedge sys_clk) begin
	memdat_16 <= mem_grain0_1[ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram1_we[0])
		mem_grain0_1[ethmac_sram1_adr1] <= ethmac_sram1_dat_w[7:0];
	memadr_53 <= ethmac_sram1_adr1;
end

assign ethmac_reader_memory1_dat_r[7:0] = memdat_16;
assign ethmac_sram1_dat_r1[7:0] = mem_grain0_1[memadr_53];

reg [7:0] mem_grain1_1[0:381];
reg [7:0] memdat_17;
reg [8:0] memadr_54;
always @(posedge sys_clk) begin
	memdat_17 <= mem_grain1_1[ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram1_we[1])
		mem_grain1_1[ethmac_sram1_adr1] <= ethmac_sram1_dat_w[15:8];
	memadr_54 <= ethmac_sram1_adr1;
end

assign ethmac_reader_memory1_dat_r[15:8] = memdat_17;
assign ethmac_sram1_dat_r1[15:8] = mem_grain1_1[memadr_54];

reg [7:0] mem_grain2_1[0:381];
reg [7:0] memdat_18;
reg [8:0] memadr_55;
always @(posedge sys_clk) begin
	memdat_18 <= mem_grain2_1[ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram1_we[2])
		mem_grain2_1[ethmac_sram1_adr1] <= ethmac_sram1_dat_w[23:16];
	memadr_55 <= ethmac_sram1_adr1;
end

assign ethmac_reader_memory1_dat_r[23:16] = memdat_18;
assign ethmac_sram1_dat_r1[23:16] = mem_grain2_1[memadr_55];

reg [7:0] mem_grain3_1[0:381];
reg [7:0] memdat_19;
reg [8:0] memadr_56;
always @(posedge sys_clk) begin
	memdat_19 <= mem_grain3_1[ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (ethmac_sram1_we[3])
		mem_grain3_1[ethmac_sram1_adr1] <= ethmac_sram1_dat_w[31:24];
	memadr_56 <= ethmac_sram1_adr1;
end

assign ethmac_reader_memory1_dat_r[31:24] = memdat_19;
assign ethmac_sram1_dat_r1[31:24] = mem_grain3_1[memadr_56];

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl0),
	.Q(xilinxasyncresetsynchronizerimpl0_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl0),
	.Q(sys_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl1),
	.Q(xilinxasyncresetsynchronizerimpl1_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl1),
	.Q(clk200_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(clk100_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl2),
	.Q(xilinxasyncresetsynchronizerimpl2_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(clk100_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl2),
	.Q(clk100_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(ethphy_reset0),
	.Q(xilinxasyncresetsynchronizerimpl3_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(ethphy_reset0),
	.Q(eth_tx_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_8 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(ethphy_reset0),
	.Q(xilinxasyncresetsynchronizerimpl4_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_9 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl4_rst_meta),
	.PRE(ethphy_reset0),
	.Q(eth_rx_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_10 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl5),
	.Q(xilinxasyncresetsynchronizerimpl5_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_11 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl5_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl5),
	.Q(hdmi_in0_pix_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_12 (
	.C(pix1p25x_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl6),
	.Q(xilinxasyncresetsynchronizerimpl6_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_13 (
	.C(pix1p25x_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl6_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl6),
	.Q(pix1p25x_rst)
);

endmodule
