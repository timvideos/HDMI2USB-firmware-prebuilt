/* Machine-generated using Migen */
module top(
	input serial_rx,
	output reg serial_tx,
	input clk100,
	input cpu_reset,
	output ddram_clock_p,
	output ddram_clock_n,
	output reg spiflash4x_cs_n,
	output reg spiflash4x_clk,
	inout [3:0] spiflash4x_dq,
	output reg ddram_cke,
	output reg ddram_ras_n,
	output reg ddram_cas_n,
	output reg ddram_we_n,
	output reg [2:0] ddram_ba,
	output reg [12:0] ddram_a,
	inout [15:0] ddram_dq,
	output [1:0] ddram_dqs,
	output [1:0] ddram_dqs_n,
	output [1:0] ddram_dm,
	output reg ddram_odt,
	input hdmi_in0_clk_p,
	input hdmi_in0_clk_n,
	input hdmi_in0_data0_p,
	input hdmi_in0_data0_n,
	input hdmi_in0_data1_p,
	input hdmi_in0_data1_n,
	input hdmi_in0_data2_p,
	input hdmi_in0_data2_n,
	input hdmi_in0_scl,
	inout hdmi_in0_sda,
	input hdmi_in1_clk_p,
	input hdmi_in1_clk_n,
	input hdmi_in1_data0_p,
	input hdmi_in1_data0_n,
	input hdmi_in1_data1_p,
	input hdmi_in1_data1_n,
	input hdmi_in1_data2_p,
	input hdmi_in1_data2_n,
	input hdmi_in1_scl,
	inout hdmi_in1_sda,
	output hdmi_out0_clk_p,
	output hdmi_out0_clk_n,
	output hdmi_out0_data0_p,
	output hdmi_out0_data0_n,
	output hdmi_out0_data1_p,
	output hdmi_out0_data1_n,
	output hdmi_out0_data2_p,
	output hdmi_out0_data2_n,
	input hdmi_out0_scl,
	input hdmi_out0_sda,
	output hdmi_out1_clk_p,
	output hdmi_out1_clk_n,
	output hdmi_out1_data0_p,
	output hdmi_out1_data0_n,
	output hdmi_out1_data1_p,
	output hdmi_out1_data1_n,
	output hdmi_out1_data2_p,
	output hdmi_out1_data2_n,
	input fx2_ifclk,
	inout [7:0] fx2_data,
	output [1:0] fx2_addr,
	input fx2_flaga,
	input fx2_flagb,
	input fx2_flagc,
	output fx2_rd_n,
	output fx2_wr_n,
	output fx2_oe_n,
	output fx2_cs_n,
	output fx2_pktend_n
);

wire [29:0] hdmi2usbsoc_hdmi2usbsoc_ibus_adr;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_ibus_dat_w;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_ibus_dat_r;
wire [3:0] hdmi2usbsoc_hdmi2usbsoc_ibus_sel;
wire hdmi2usbsoc_hdmi2usbsoc_ibus_cyc;
wire hdmi2usbsoc_hdmi2usbsoc_ibus_stb;
wire hdmi2usbsoc_hdmi2usbsoc_ibus_ack;
wire hdmi2usbsoc_hdmi2usbsoc_ibus_we;
wire [2:0] hdmi2usbsoc_hdmi2usbsoc_ibus_cti;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_ibus_bte;
wire hdmi2usbsoc_hdmi2usbsoc_ibus_err;
wire [29:0] hdmi2usbsoc_hdmi2usbsoc_dbus_adr;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_dbus_dat_w;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_dbus_dat_r;
wire [3:0] hdmi2usbsoc_hdmi2usbsoc_dbus_sel;
wire hdmi2usbsoc_hdmi2usbsoc_dbus_cyc;
wire hdmi2usbsoc_hdmi2usbsoc_dbus_stb;
wire hdmi2usbsoc_hdmi2usbsoc_dbus_ack;
wire hdmi2usbsoc_hdmi2usbsoc_dbus_we;
wire [2:0] hdmi2usbsoc_hdmi2usbsoc_dbus_cti;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_dbus_bte;
wire hdmi2usbsoc_hdmi2usbsoc_dbus_err;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_interrupt = 32'd0;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_i_adr_o;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_d_adr_o;
wire [29:0] hdmi2usbsoc_hdmi2usbsoc_rom_bus_adr;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_rom_bus_dat_w;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_rom_bus_dat_r;
wire [3:0] hdmi2usbsoc_hdmi2usbsoc_rom_bus_sel;
wire hdmi2usbsoc_hdmi2usbsoc_rom_bus_cyc;
wire hdmi2usbsoc_hdmi2usbsoc_rom_bus_stb;
reg hdmi2usbsoc_hdmi2usbsoc_rom_bus_ack = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_rom_bus_we;
wire [2:0] hdmi2usbsoc_hdmi2usbsoc_rom_bus_cti;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_rom_bus_bte;
reg hdmi2usbsoc_hdmi2usbsoc_rom_bus_err = 1'd0;
wire [12:0] hdmi2usbsoc_hdmi2usbsoc_rom_adr;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_rom_dat_r;
wire [29:0] hdmi2usbsoc_hdmi2usbsoc_sram_bus_adr;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_sram_bus_dat_w;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_sram_bus_dat_r;
wire [3:0] hdmi2usbsoc_hdmi2usbsoc_sram_bus_sel;
wire hdmi2usbsoc_hdmi2usbsoc_sram_bus_cyc;
wire hdmi2usbsoc_hdmi2usbsoc_sram_bus_stb;
reg hdmi2usbsoc_hdmi2usbsoc_sram_bus_ack = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_sram_bus_we;
wire [2:0] hdmi2usbsoc_hdmi2usbsoc_sram_bus_cti;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_sram_bus_bte;
reg hdmi2usbsoc_hdmi2usbsoc_sram_bus_err = 1'd0;
wire [11:0] hdmi2usbsoc_hdmi2usbsoc_sram_adr;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_sram_dat_r;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_sram_we = 4'd0;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_sram_dat_w;
reg [13:0] hdmi2usbsoc_hdmi2usbsoc_interface_adr = 14'd0;
reg hdmi2usbsoc_hdmi2usbsoc_interface_we = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi2usbsoc_interface_dat_w = 8'd0;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_interface_dat_r;
wire [29:0] hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_adr;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_dat_w;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_dat_r = 32'd0;
wire [3:0] hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_sel;
wire hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_cyc;
wire hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_stb;
reg hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_ack = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_we;
wire [2:0] hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_cti;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_bte;
reg hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_err = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi2usbsoc_counter = 2'd0;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full = 32'd6597069;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_re = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_valid;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_ready = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_last;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_payload_data;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_reg = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_bitcount = 4'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_busy = 1'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_valid = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_ready;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_first = 1'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_last = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_payload_data = 8'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_rx = 32'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_r = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_reg = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_bitcount = 4'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_busy = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_re;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_r;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_w;
wire hdmi2usbsoc_hdmi2usbsoc_uart_txfull_status;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rxempty_status;
wire hdmi2usbsoc_hdmi2usbsoc_uart_irq;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_status;
reg hdmi2usbsoc_hdmi2usbsoc_uart_tx_pending = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_trigger;
reg hdmi2usbsoc_hdmi2usbsoc_uart_tx_clear = 1'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_tx_old_trigger = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_status;
reg hdmi2usbsoc_hdmi2usbsoc_uart_rx_pending = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_trigger;
reg hdmi2usbsoc_hdmi2usbsoc_uart_rx_clear = 1'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_rx_old_trigger = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_status_re;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_uart_status_r;
reg [1:0] hdmi2usbsoc_hdmi2usbsoc_uart_status_w = 2'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_pending_re;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_uart_pending_r;
reg [1:0] hdmi2usbsoc_hdmi2usbsoc_uart_pending_w = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi2usbsoc_uart_storage_full = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi2usbsoc_uart_storage;
reg hdmi2usbsoc_hdmi2usbsoc_uart_re = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_valid;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_ready;
reg hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_last = 1'd0;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_valid;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_ready;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_dout;
reg [4:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level = 5'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_replace = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_produce = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_consume = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_adr = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_do_read;
wire [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_last;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_valid;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_ready;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_last;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_valid;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_ready;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_dout;
reg [4:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level = 5'd0;
reg hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_replace = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_produce = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_consume = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_adr = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_do_read;
wire [3:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_last;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_load_re = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_reload_re = 1'd0;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_en_re = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_update_value_re;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_update_value_r;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_update_value_w = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_timer0_value_status = 32'd0;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_irq;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_zero_status;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_zero_pending = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_zero_trigger;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_zero_clear = 1'd0;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_zero_old_trigger = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_status_re;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_status_r;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_status_w;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_re;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_r;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_w;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage;
reg hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_re = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi2usbsoc_timer0_value = 32'd0;
wire [29:0] hdmi2usbsoc_interface0_wb_sdram_adr;
wire [31:0] hdmi2usbsoc_interface0_wb_sdram_dat_w;
reg [31:0] hdmi2usbsoc_interface0_wb_sdram_dat_r = 32'd0;
wire [3:0] hdmi2usbsoc_interface0_wb_sdram_sel;
wire hdmi2usbsoc_interface0_wb_sdram_cyc;
wire hdmi2usbsoc_interface0_wb_sdram_stb;
reg hdmi2usbsoc_interface0_wb_sdram_ack = 1'd0;
wire hdmi2usbsoc_interface0_wb_sdram_we;
wire [2:0] hdmi2usbsoc_interface0_wb_sdram_cti;
wire [1:0] hdmi2usbsoc_interface0_wb_sdram_bte;
reg hdmi2usbsoc_interface0_wb_sdram_err = 1'd0;
wire sys_clk;
wire sys_rst;
wire sdram_half_clk;
reg sdram_half_rst = 1'd0;
wire sdram_full_wr_clk;
wire sdram_full_rd_clk;
wire base50_clk;
wire base50_rst;
(* keep = "true" *) wire encoder_clk;
wire encoder_rst;
reg hdmi2usbsoc_crg_reset = 1'd0;
wire hdmi2usbsoc_crg_clk100a;
wire hdmi2usbsoc_crg_clk100b;
wire hdmi2usbsoc_crg_unbuf_sdram_full;
wire hdmi2usbsoc_crg_unbuf_sdram_half_a;
wire hdmi2usbsoc_crg_unbuf_sdram_half_b;
wire hdmi2usbsoc_crg_unbuf_encoder;
wire hdmi2usbsoc_crg_unbuf_sys;
wire hdmi2usbsoc_crg_unbuf_unused;
wire hdmi2usbsoc_crg_pll_lckd;
wire hdmi2usbsoc_crg_pll_fb;
wire por_clk;
wire por_rst;
reg [10:0] hdmi2usbsoc_crg_por = 11'd2047;
wire hdmi2usbsoc_crg_clk4x_wr_strb;
wire hdmi2usbsoc_crg_clk4x_rd_strb;
wire hdmi2usbsoc_crg_clk_sdram_half_shifted;
wire hdmi2usbsoc_crg_output_clk;
wire hdmi2usbsoc_crg_dcm_base50_locked;
reg [56:0] hdmi2usbsoc_dna_status = 57'd0;
wire hdmi2usbsoc_dna_do;
reg [6:0] hdmi2usbsoc_dna_cnt = 7'd0;
wire [159:0] hdmi2usbsoc_git_status;
wire [63:0] hdmi2usbsoc_platform_status;
wire [63:0] hdmi2usbsoc_target_status;
wire [29:0] hdmi2usbsoc_bus_adr;
wire [31:0] hdmi2usbsoc_bus_dat_w;
wire [31:0] hdmi2usbsoc_bus_dat_r;
wire [3:0] hdmi2usbsoc_bus_sel;
wire hdmi2usbsoc_bus_cyc;
wire hdmi2usbsoc_bus_stb;
reg hdmi2usbsoc_bus_ack = 1'd0;
wire hdmi2usbsoc_bus_we;
wire [2:0] hdmi2usbsoc_bus_cti;
wire [1:0] hdmi2usbsoc_bus_bte;
reg hdmi2usbsoc_bus_err = 1'd0;
reg [3:0] hdmi2usbsoc_bitbang_storage_full = 4'd0;
wire [3:0] hdmi2usbsoc_bitbang_storage;
reg hdmi2usbsoc_bitbang_re = 1'd0;
reg hdmi2usbsoc_status = 1'd0;
reg hdmi2usbsoc_bitbang_en_storage_full = 1'd0;
wire hdmi2usbsoc_bitbang_en_storage;
reg hdmi2usbsoc_bitbang_en_re = 1'd0;
reg hdmi2usbsoc_cs_n = 1'd1;
reg hdmi2usbsoc_clk = 1'd0;
reg hdmi2usbsoc_dq_oe = 1'd0;
reg [3:0] hdmi2usbsoc_o = 4'd0;
reg hdmi2usbsoc_oe = 1'd0;
wire [3:0] hdmi2usbsoc_i0;
reg [31:0] hdmi2usbsoc_sr = 32'd0;
reg [1:0] hdmi2usbsoc_i1 = 2'd0;
reg [3:0] hdmi2usbsoc_dqi = 4'd0;
reg [7:0] hdmi2usbsoc_counter = 8'd0;
wire [12:0] hdmi2usbsoc_ddrphy_dfi_p0_address;
wire [2:0] hdmi2usbsoc_ddrphy_dfi_p0_bank;
wire hdmi2usbsoc_ddrphy_dfi_p0_cas_n;
wire hdmi2usbsoc_ddrphy_dfi_p0_cs_n;
wire hdmi2usbsoc_ddrphy_dfi_p0_ras_n;
wire hdmi2usbsoc_ddrphy_dfi_p0_we_n;
wire hdmi2usbsoc_ddrphy_dfi_p0_cke;
wire hdmi2usbsoc_ddrphy_dfi_p0_odt;
wire hdmi2usbsoc_ddrphy_dfi_p0_reset_n;
wire [31:0] hdmi2usbsoc_ddrphy_dfi_p0_wrdata;
wire hdmi2usbsoc_ddrphy_dfi_p0_wrdata_en;
wire [3:0] hdmi2usbsoc_ddrphy_dfi_p0_wrdata_mask;
wire hdmi2usbsoc_ddrphy_dfi_p0_rddata_en;
wire [31:0] hdmi2usbsoc_ddrphy_dfi_p0_rddata;
wire hdmi2usbsoc_ddrphy_dfi_p0_rddata_valid;
wire [12:0] hdmi2usbsoc_ddrphy_dfi_p1_address;
wire [2:0] hdmi2usbsoc_ddrphy_dfi_p1_bank;
wire hdmi2usbsoc_ddrphy_dfi_p1_cas_n;
wire hdmi2usbsoc_ddrphy_dfi_p1_cs_n;
wire hdmi2usbsoc_ddrphy_dfi_p1_ras_n;
wire hdmi2usbsoc_ddrphy_dfi_p1_we_n;
wire hdmi2usbsoc_ddrphy_dfi_p1_cke;
wire hdmi2usbsoc_ddrphy_dfi_p1_odt;
wire hdmi2usbsoc_ddrphy_dfi_p1_reset_n;
wire [31:0] hdmi2usbsoc_ddrphy_dfi_p1_wrdata;
wire hdmi2usbsoc_ddrphy_dfi_p1_wrdata_en;
wire [3:0] hdmi2usbsoc_ddrphy_dfi_p1_wrdata_mask;
wire hdmi2usbsoc_ddrphy_dfi_p1_rddata_en;
wire [31:0] hdmi2usbsoc_ddrphy_dfi_p1_rddata;
wire hdmi2usbsoc_ddrphy_dfi_p1_rddata_valid;
wire hdmi2usbsoc_ddrphy_clk4x_wr_strb;
wire hdmi2usbsoc_ddrphy_clk4x_rd_strb;
reg hdmi2usbsoc_ddrphy_phase_sel = 1'd0;
reg hdmi2usbsoc_ddrphy_phase_half = 1'd0;
reg hdmi2usbsoc_ddrphy_phase_sys = 1'd0;
reg [12:0] hdmi2usbsoc_ddrphy_record0_address = 13'd0;
reg [2:0] hdmi2usbsoc_ddrphy_record0_bank = 3'd0;
reg hdmi2usbsoc_ddrphy_record0_cas_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record0_cs_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record0_ras_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record0_we_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record0_cke = 1'd0;
reg hdmi2usbsoc_ddrphy_record0_odt = 1'd0;
reg hdmi2usbsoc_ddrphy_record0_reset_n = 1'd0;
reg [12:0] hdmi2usbsoc_ddrphy_record1_address = 13'd0;
reg [2:0] hdmi2usbsoc_ddrphy_record1_bank = 3'd0;
reg hdmi2usbsoc_ddrphy_record1_cas_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record1_cs_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record1_ras_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record1_we_n = 1'd0;
reg hdmi2usbsoc_ddrphy_record1_cke = 1'd0;
reg hdmi2usbsoc_ddrphy_record1_odt = 1'd0;
reg hdmi2usbsoc_ddrphy_record1_reset_n = 1'd0;
reg [3:0] hdmi2usbsoc_ddrphy_bitslip_cnt = 4'd0;
reg hdmi2usbsoc_ddrphy_bitslip_inc = 1'd0;
wire hdmi2usbsoc_ddrphy_sdram_half_clk_n;
reg hdmi2usbsoc_ddrphy_postamble = 1'd0;
wire hdmi2usbsoc_ddrphy_drive_dqs;
wire hdmi2usbsoc_ddrphy_dqs_t_d0;
wire hdmi2usbsoc_ddrphy_dqs_t_d1;
wire [1:0] hdmi2usbsoc_ddrphy_dqs_o;
wire [1:0] hdmi2usbsoc_ddrphy_dqs_t;
wire [31:0] hdmi2usbsoc_ddrphy_record0_wrdata;
wire hdmi2usbsoc_ddrphy_record0_wrdata_en;
wire [3:0] hdmi2usbsoc_ddrphy_record0_wrdata_mask;
wire hdmi2usbsoc_ddrphy_record0_rddata_en;
wire [31:0] hdmi2usbsoc_ddrphy_record0_rddata;
wire [31:0] hdmi2usbsoc_ddrphy_record1_wrdata;
wire hdmi2usbsoc_ddrphy_record1_wrdata_en;
wire [3:0] hdmi2usbsoc_ddrphy_record1_wrdata_mask;
wire hdmi2usbsoc_ddrphy_record1_rddata_en;
wire [31:0] hdmi2usbsoc_ddrphy_record1_rddata;
reg [31:0] hdmi2usbsoc_ddrphy_record2_wrdata = 32'd0;
reg [3:0] hdmi2usbsoc_ddrphy_record2_wrdata_mask = 4'd0;
reg [31:0] hdmi2usbsoc_ddrphy_record3_wrdata = 32'd0;
reg [3:0] hdmi2usbsoc_ddrphy_record3_wrdata_mask = 4'd0;
wire hdmi2usbsoc_ddrphy_drive_dq;
wire hdmi2usbsoc_ddrphy_drive_dq_n0;
reg hdmi2usbsoc_ddrphy_drive_dq_n1 = 1'd0;
wire [15:0] hdmi2usbsoc_ddrphy_dq_t;
wire [15:0] hdmi2usbsoc_ddrphy_dq_o;
wire [15:0] hdmi2usbsoc_ddrphy_dq_i;
wire hdmi2usbsoc_ddrphy_wrdata_en;
reg hdmi2usbsoc_ddrphy_wrdata_en_d = 1'd0;
reg [2:0] hdmi2usbsoc_ddrphy_r_dfi_wrdata_en = 3'd0;
wire hdmi2usbsoc_ddrphy_rddata_en;
reg [4:0] hdmi2usbsoc_ddrphy_rddata_sr = 5'd0;
wire [12:0] hdmi2usbsoc_sdram_inti_p0_address;
wire [2:0] hdmi2usbsoc_sdram_inti_p0_bank;
reg hdmi2usbsoc_sdram_inti_p0_cas_n = 1'd1;
reg hdmi2usbsoc_sdram_inti_p0_cs_n = 1'd1;
reg hdmi2usbsoc_sdram_inti_p0_ras_n = 1'd1;
reg hdmi2usbsoc_sdram_inti_p0_we_n = 1'd1;
wire hdmi2usbsoc_sdram_inti_p0_cke;
wire hdmi2usbsoc_sdram_inti_p0_odt;
wire hdmi2usbsoc_sdram_inti_p0_reset_n;
wire [31:0] hdmi2usbsoc_sdram_inti_p0_wrdata;
wire hdmi2usbsoc_sdram_inti_p0_wrdata_en;
wire [3:0] hdmi2usbsoc_sdram_inti_p0_wrdata_mask;
wire hdmi2usbsoc_sdram_inti_p0_rddata_en;
reg [31:0] hdmi2usbsoc_sdram_inti_p0_rddata = 32'd0;
reg hdmi2usbsoc_sdram_inti_p0_rddata_valid = 1'd0;
wire [12:0] hdmi2usbsoc_sdram_inti_p1_address;
wire [2:0] hdmi2usbsoc_sdram_inti_p1_bank;
reg hdmi2usbsoc_sdram_inti_p1_cas_n = 1'd1;
reg hdmi2usbsoc_sdram_inti_p1_cs_n = 1'd1;
reg hdmi2usbsoc_sdram_inti_p1_ras_n = 1'd1;
reg hdmi2usbsoc_sdram_inti_p1_we_n = 1'd1;
wire hdmi2usbsoc_sdram_inti_p1_cke;
wire hdmi2usbsoc_sdram_inti_p1_odt;
wire hdmi2usbsoc_sdram_inti_p1_reset_n;
wire [31:0] hdmi2usbsoc_sdram_inti_p1_wrdata;
wire hdmi2usbsoc_sdram_inti_p1_wrdata_en;
wire [3:0] hdmi2usbsoc_sdram_inti_p1_wrdata_mask;
wire hdmi2usbsoc_sdram_inti_p1_rddata_en;
reg [31:0] hdmi2usbsoc_sdram_inti_p1_rddata = 32'd0;
reg hdmi2usbsoc_sdram_inti_p1_rddata_valid = 1'd0;
wire [12:0] hdmi2usbsoc_sdram_slave_p0_address;
wire [2:0] hdmi2usbsoc_sdram_slave_p0_bank;
wire hdmi2usbsoc_sdram_slave_p0_cas_n;
wire hdmi2usbsoc_sdram_slave_p0_cs_n;
wire hdmi2usbsoc_sdram_slave_p0_ras_n;
wire hdmi2usbsoc_sdram_slave_p0_we_n;
wire hdmi2usbsoc_sdram_slave_p0_cke;
wire hdmi2usbsoc_sdram_slave_p0_odt;
wire hdmi2usbsoc_sdram_slave_p0_reset_n;
wire [31:0] hdmi2usbsoc_sdram_slave_p0_wrdata;
wire hdmi2usbsoc_sdram_slave_p0_wrdata_en;
wire [3:0] hdmi2usbsoc_sdram_slave_p0_wrdata_mask;
wire hdmi2usbsoc_sdram_slave_p0_rddata_en;
reg [31:0] hdmi2usbsoc_sdram_slave_p0_rddata = 32'd0;
reg hdmi2usbsoc_sdram_slave_p0_rddata_valid = 1'd0;
wire [12:0] hdmi2usbsoc_sdram_slave_p1_address;
wire [2:0] hdmi2usbsoc_sdram_slave_p1_bank;
wire hdmi2usbsoc_sdram_slave_p1_cas_n;
wire hdmi2usbsoc_sdram_slave_p1_cs_n;
wire hdmi2usbsoc_sdram_slave_p1_ras_n;
wire hdmi2usbsoc_sdram_slave_p1_we_n;
wire hdmi2usbsoc_sdram_slave_p1_cke;
wire hdmi2usbsoc_sdram_slave_p1_odt;
wire hdmi2usbsoc_sdram_slave_p1_reset_n;
wire [31:0] hdmi2usbsoc_sdram_slave_p1_wrdata;
wire hdmi2usbsoc_sdram_slave_p1_wrdata_en;
wire [3:0] hdmi2usbsoc_sdram_slave_p1_wrdata_mask;
wire hdmi2usbsoc_sdram_slave_p1_rddata_en;
reg [31:0] hdmi2usbsoc_sdram_slave_p1_rddata = 32'd0;
reg hdmi2usbsoc_sdram_slave_p1_rddata_valid = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_master_p0_address = 13'd0;
reg [2:0] hdmi2usbsoc_sdram_master_p0_bank = 3'd0;
reg hdmi2usbsoc_sdram_master_p0_cas_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p0_cs_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p0_ras_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p0_we_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p0_cke = 1'd0;
reg hdmi2usbsoc_sdram_master_p0_odt = 1'd0;
reg hdmi2usbsoc_sdram_master_p0_reset_n = 1'd0;
reg [31:0] hdmi2usbsoc_sdram_master_p0_wrdata = 32'd0;
reg hdmi2usbsoc_sdram_master_p0_wrdata_en = 1'd0;
reg [3:0] hdmi2usbsoc_sdram_master_p0_wrdata_mask = 4'd0;
reg hdmi2usbsoc_sdram_master_p0_rddata_en = 1'd0;
wire [31:0] hdmi2usbsoc_sdram_master_p0_rddata;
wire hdmi2usbsoc_sdram_master_p0_rddata_valid;
reg [12:0] hdmi2usbsoc_sdram_master_p1_address = 13'd0;
reg [2:0] hdmi2usbsoc_sdram_master_p1_bank = 3'd0;
reg hdmi2usbsoc_sdram_master_p1_cas_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p1_cs_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p1_ras_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p1_we_n = 1'd1;
reg hdmi2usbsoc_sdram_master_p1_cke = 1'd0;
reg hdmi2usbsoc_sdram_master_p1_odt = 1'd0;
reg hdmi2usbsoc_sdram_master_p1_reset_n = 1'd0;
reg [31:0] hdmi2usbsoc_sdram_master_p1_wrdata = 32'd0;
reg hdmi2usbsoc_sdram_master_p1_wrdata_en = 1'd0;
reg [3:0] hdmi2usbsoc_sdram_master_p1_wrdata_mask = 4'd0;
reg hdmi2usbsoc_sdram_master_p1_rddata_en = 1'd0;
wire [31:0] hdmi2usbsoc_sdram_master_p1_rddata;
wire hdmi2usbsoc_sdram_master_p1_rddata_valid;
reg [3:0] hdmi2usbsoc_sdram_storage_full = 4'd0;
wire [3:0] hdmi2usbsoc_sdram_storage;
reg hdmi2usbsoc_sdram_re = 1'd0;
reg [5:0] hdmi2usbsoc_sdram_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] hdmi2usbsoc_sdram_phaseinjector0_command_storage;
reg hdmi2usbsoc_sdram_phaseinjector0_command_re = 1'd0;
wire hdmi2usbsoc_sdram_phaseinjector0_command_issue_re;
wire hdmi2usbsoc_sdram_phaseinjector0_command_issue_r;
reg hdmi2usbsoc_sdram_phaseinjector0_command_issue_w = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_phaseinjector0_address_storage_full = 13'd0;
wire [12:0] hdmi2usbsoc_sdram_phaseinjector0_address_storage;
reg hdmi2usbsoc_sdram_phaseinjector0_address_re = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] hdmi2usbsoc_sdram_phaseinjector0_baddress_storage;
reg hdmi2usbsoc_sdram_phaseinjector0_baddress_re = 1'd0;
reg [31:0] hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage;
reg hdmi2usbsoc_sdram_phaseinjector0_wrdata_re = 1'd0;
reg [31:0] hdmi2usbsoc_sdram_phaseinjector0_status = 32'd0;
reg [5:0] hdmi2usbsoc_sdram_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] hdmi2usbsoc_sdram_phaseinjector1_command_storage;
reg hdmi2usbsoc_sdram_phaseinjector1_command_re = 1'd0;
wire hdmi2usbsoc_sdram_phaseinjector1_command_issue_re;
wire hdmi2usbsoc_sdram_phaseinjector1_command_issue_r;
reg hdmi2usbsoc_sdram_phaseinjector1_command_issue_w = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_phaseinjector1_address_storage_full = 13'd0;
wire [12:0] hdmi2usbsoc_sdram_phaseinjector1_address_storage;
reg hdmi2usbsoc_sdram_phaseinjector1_address_re = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] hdmi2usbsoc_sdram_phaseinjector1_baddress_storage;
reg hdmi2usbsoc_sdram_phaseinjector1_baddress_re = 1'd0;
reg [31:0] hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage;
reg hdmi2usbsoc_sdram_phaseinjector1_wrdata_re = 1'd0;
reg [31:0] hdmi2usbsoc_sdram_phaseinjector1_status = 32'd0;
reg [12:0] hdmi2usbsoc_sdram_dfi_p0_address = 13'd0;
reg [2:0] hdmi2usbsoc_sdram_dfi_p0_bank = 3'd0;
reg hdmi2usbsoc_sdram_dfi_p0_cas_n = 1'd1;
wire hdmi2usbsoc_sdram_dfi_p0_cs_n;
reg hdmi2usbsoc_sdram_dfi_p0_ras_n = 1'd1;
reg hdmi2usbsoc_sdram_dfi_p0_we_n = 1'd1;
wire hdmi2usbsoc_sdram_dfi_p0_cke;
wire hdmi2usbsoc_sdram_dfi_p0_odt;
wire hdmi2usbsoc_sdram_dfi_p0_reset_n;
wire [31:0] hdmi2usbsoc_sdram_dfi_p0_wrdata;
reg hdmi2usbsoc_sdram_dfi_p0_wrdata_en = 1'd0;
wire [3:0] hdmi2usbsoc_sdram_dfi_p0_wrdata_mask;
reg hdmi2usbsoc_sdram_dfi_p0_rddata_en = 1'd0;
wire [31:0] hdmi2usbsoc_sdram_dfi_p0_rddata;
wire hdmi2usbsoc_sdram_dfi_p0_rddata_valid;
reg [12:0] hdmi2usbsoc_sdram_dfi_p1_address = 13'd0;
reg [2:0] hdmi2usbsoc_sdram_dfi_p1_bank = 3'd0;
reg hdmi2usbsoc_sdram_dfi_p1_cas_n = 1'd1;
wire hdmi2usbsoc_sdram_dfi_p1_cs_n;
reg hdmi2usbsoc_sdram_dfi_p1_ras_n = 1'd1;
reg hdmi2usbsoc_sdram_dfi_p1_we_n = 1'd1;
wire hdmi2usbsoc_sdram_dfi_p1_cke;
wire hdmi2usbsoc_sdram_dfi_p1_odt;
wire hdmi2usbsoc_sdram_dfi_p1_reset_n;
wire [31:0] hdmi2usbsoc_sdram_dfi_p1_wrdata;
reg hdmi2usbsoc_sdram_dfi_p1_wrdata_en = 1'd0;
wire [3:0] hdmi2usbsoc_sdram_dfi_p1_wrdata_mask;
reg hdmi2usbsoc_sdram_dfi_p1_rddata_en = 1'd0;
wire [31:0] hdmi2usbsoc_sdram_dfi_p1_rddata;
wire hdmi2usbsoc_sdram_dfi_p1_rddata_valid;
wire hdmi2usbsoc_sdram_interface_bank0_valid;
wire hdmi2usbsoc_sdram_interface_bank0_ready;
wire hdmi2usbsoc_sdram_interface_bank0_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank0_adr;
wire hdmi2usbsoc_sdram_interface_bank0_lock;
wire hdmi2usbsoc_sdram_interface_bank0_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank0_rdata_valid;
wire hdmi2usbsoc_sdram_interface_bank1_valid;
wire hdmi2usbsoc_sdram_interface_bank1_ready;
wire hdmi2usbsoc_sdram_interface_bank1_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank1_adr;
wire hdmi2usbsoc_sdram_interface_bank1_lock;
wire hdmi2usbsoc_sdram_interface_bank1_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank1_rdata_valid;
wire hdmi2usbsoc_sdram_interface_bank2_valid;
wire hdmi2usbsoc_sdram_interface_bank2_ready;
wire hdmi2usbsoc_sdram_interface_bank2_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank2_adr;
wire hdmi2usbsoc_sdram_interface_bank2_lock;
wire hdmi2usbsoc_sdram_interface_bank2_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank2_rdata_valid;
wire hdmi2usbsoc_sdram_interface_bank3_valid;
wire hdmi2usbsoc_sdram_interface_bank3_ready;
wire hdmi2usbsoc_sdram_interface_bank3_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank3_adr;
wire hdmi2usbsoc_sdram_interface_bank3_lock;
wire hdmi2usbsoc_sdram_interface_bank3_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank3_rdata_valid;
wire hdmi2usbsoc_sdram_interface_bank4_valid;
wire hdmi2usbsoc_sdram_interface_bank4_ready;
wire hdmi2usbsoc_sdram_interface_bank4_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank4_adr;
wire hdmi2usbsoc_sdram_interface_bank4_lock;
wire hdmi2usbsoc_sdram_interface_bank4_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank4_rdata_valid;
wire hdmi2usbsoc_sdram_interface_bank5_valid;
wire hdmi2usbsoc_sdram_interface_bank5_ready;
wire hdmi2usbsoc_sdram_interface_bank5_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank5_adr;
wire hdmi2usbsoc_sdram_interface_bank5_lock;
wire hdmi2usbsoc_sdram_interface_bank5_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank5_rdata_valid;
wire hdmi2usbsoc_sdram_interface_bank6_valid;
wire hdmi2usbsoc_sdram_interface_bank6_ready;
wire hdmi2usbsoc_sdram_interface_bank6_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank6_adr;
wire hdmi2usbsoc_sdram_interface_bank6_lock;
wire hdmi2usbsoc_sdram_interface_bank6_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank6_rdata_valid;
wire hdmi2usbsoc_sdram_interface_bank7_valid;
wire hdmi2usbsoc_sdram_interface_bank7_ready;
wire hdmi2usbsoc_sdram_interface_bank7_we;
wire [20:0] hdmi2usbsoc_sdram_interface_bank7_adr;
wire hdmi2usbsoc_sdram_interface_bank7_lock;
wire hdmi2usbsoc_sdram_interface_bank7_wdata_ready;
wire hdmi2usbsoc_sdram_interface_bank7_rdata_valid;
reg [63:0] hdmi2usbsoc_sdram_interface_wdata = 64'd0;
reg [7:0] hdmi2usbsoc_sdram_interface_wdata_we = 8'd0;
wire [63:0] hdmi2usbsoc_sdram_interface_rdata;
reg hdmi2usbsoc_sdram_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_cmd_ready = 1'd0;
reg hdmi2usbsoc_sdram_cmd_last = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_cmd_payload_a = 13'd0;
reg [2:0] hdmi2usbsoc_sdram_cmd_payload_ba = 3'd0;
reg hdmi2usbsoc_sdram_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_cmd_payload_is_write = 1'd0;
reg hdmi2usbsoc_sdram_seq_start = 1'd0;
reg hdmi2usbsoc_sdram_seq_done = 1'd0;
reg [3:0] hdmi2usbsoc_sdram_counter = 4'd0;
wire hdmi2usbsoc_sdram_wait;
wire hdmi2usbsoc_sdram_done;
reg [9:0] hdmi2usbsoc_sdram_count = 10'd585;
wire hdmi2usbsoc_sdram_bankmachine0_req_valid;
wire hdmi2usbsoc_sdram_bankmachine0_req_ready;
wire hdmi2usbsoc_sdram_bankmachine0_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine0_req_adr;
wire hdmi2usbsoc_sdram_bankmachine0_req_lock;
reg hdmi2usbsoc_sdram_bankmachine0_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine0_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine0_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine0_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine0_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine0_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine0_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine0_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine0_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine0_source_valid;
wire hdmi2usbsoc_sdram_bankmachine0_source_ready;
wire hdmi2usbsoc_sdram_bankmachine0_source_first;
wire hdmi2usbsoc_sdram_bankmachine0_source_last;
wire hdmi2usbsoc_sdram_bankmachine0_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine0_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine0_syncfifo0_we;
wire hdmi2usbsoc_sdram_bankmachine0_syncfifo0_writable;
wire hdmi2usbsoc_sdram_bankmachine0_syncfifo0_re;
wire hdmi2usbsoc_sdram_bankmachine0_syncfifo0_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine0_syncfifo0_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine0_syncfifo0_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine0_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine0_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine0_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine0_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine0_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine0_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine0_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine0_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine0_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine0_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine0_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine0_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine0_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine0_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine0_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine0_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine0_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine0_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine0_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine0_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine0_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine0_hit;
reg hdmi2usbsoc_sdram_bankmachine0_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine0_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine0_wait;
wire hdmi2usbsoc_sdram_bankmachine0_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine0_count = 3'd4;
wire hdmi2usbsoc_sdram_bankmachine1_req_valid;
wire hdmi2usbsoc_sdram_bankmachine1_req_ready;
wire hdmi2usbsoc_sdram_bankmachine1_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine1_req_adr;
wire hdmi2usbsoc_sdram_bankmachine1_req_lock;
reg hdmi2usbsoc_sdram_bankmachine1_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine1_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine1_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine1_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine1_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine1_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine1_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine1_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine1_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine1_source_valid;
wire hdmi2usbsoc_sdram_bankmachine1_source_ready;
wire hdmi2usbsoc_sdram_bankmachine1_source_first;
wire hdmi2usbsoc_sdram_bankmachine1_source_last;
wire hdmi2usbsoc_sdram_bankmachine1_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine1_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine1_syncfifo1_we;
wire hdmi2usbsoc_sdram_bankmachine1_syncfifo1_writable;
wire hdmi2usbsoc_sdram_bankmachine1_syncfifo1_re;
wire hdmi2usbsoc_sdram_bankmachine1_syncfifo1_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine1_syncfifo1_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine1_syncfifo1_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine1_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine1_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine1_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine1_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine1_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine1_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine1_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine1_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine1_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine1_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine1_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine1_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine1_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine1_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine1_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine1_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine1_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine1_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine1_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine1_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine1_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine1_hit;
reg hdmi2usbsoc_sdram_bankmachine1_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine1_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine1_wait;
wire hdmi2usbsoc_sdram_bankmachine1_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine1_count = 3'd4;
wire hdmi2usbsoc_sdram_bankmachine2_req_valid;
wire hdmi2usbsoc_sdram_bankmachine2_req_ready;
wire hdmi2usbsoc_sdram_bankmachine2_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine2_req_adr;
wire hdmi2usbsoc_sdram_bankmachine2_req_lock;
reg hdmi2usbsoc_sdram_bankmachine2_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine2_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine2_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine2_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine2_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine2_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine2_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine2_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine2_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine2_source_valid;
wire hdmi2usbsoc_sdram_bankmachine2_source_ready;
wire hdmi2usbsoc_sdram_bankmachine2_source_first;
wire hdmi2usbsoc_sdram_bankmachine2_source_last;
wire hdmi2usbsoc_sdram_bankmachine2_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine2_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine2_syncfifo2_we;
wire hdmi2usbsoc_sdram_bankmachine2_syncfifo2_writable;
wire hdmi2usbsoc_sdram_bankmachine2_syncfifo2_re;
wire hdmi2usbsoc_sdram_bankmachine2_syncfifo2_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine2_syncfifo2_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine2_syncfifo2_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine2_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine2_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine2_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine2_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine2_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine2_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine2_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine2_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine2_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine2_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine2_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine2_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine2_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine2_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine2_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine2_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine2_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine2_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine2_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine2_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine2_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine2_hit;
reg hdmi2usbsoc_sdram_bankmachine2_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine2_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine2_wait;
wire hdmi2usbsoc_sdram_bankmachine2_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine2_count = 3'd4;
wire hdmi2usbsoc_sdram_bankmachine3_req_valid;
wire hdmi2usbsoc_sdram_bankmachine3_req_ready;
wire hdmi2usbsoc_sdram_bankmachine3_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine3_req_adr;
wire hdmi2usbsoc_sdram_bankmachine3_req_lock;
reg hdmi2usbsoc_sdram_bankmachine3_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine3_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine3_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine3_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine3_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine3_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine3_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine3_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine3_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine3_source_valid;
wire hdmi2usbsoc_sdram_bankmachine3_source_ready;
wire hdmi2usbsoc_sdram_bankmachine3_source_first;
wire hdmi2usbsoc_sdram_bankmachine3_source_last;
wire hdmi2usbsoc_sdram_bankmachine3_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine3_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine3_syncfifo3_we;
wire hdmi2usbsoc_sdram_bankmachine3_syncfifo3_writable;
wire hdmi2usbsoc_sdram_bankmachine3_syncfifo3_re;
wire hdmi2usbsoc_sdram_bankmachine3_syncfifo3_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine3_syncfifo3_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine3_syncfifo3_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine3_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine3_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine3_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine3_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine3_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine3_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine3_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine3_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine3_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine3_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine3_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine3_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine3_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine3_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine3_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine3_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine3_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine3_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine3_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine3_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine3_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine3_hit;
reg hdmi2usbsoc_sdram_bankmachine3_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine3_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine3_wait;
wire hdmi2usbsoc_sdram_bankmachine3_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine3_count = 3'd4;
wire hdmi2usbsoc_sdram_bankmachine4_req_valid;
wire hdmi2usbsoc_sdram_bankmachine4_req_ready;
wire hdmi2usbsoc_sdram_bankmachine4_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine4_req_adr;
wire hdmi2usbsoc_sdram_bankmachine4_req_lock;
reg hdmi2usbsoc_sdram_bankmachine4_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine4_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine4_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine4_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine4_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine4_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine4_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine4_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine4_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine4_source_valid;
wire hdmi2usbsoc_sdram_bankmachine4_source_ready;
wire hdmi2usbsoc_sdram_bankmachine4_source_first;
wire hdmi2usbsoc_sdram_bankmachine4_source_last;
wire hdmi2usbsoc_sdram_bankmachine4_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine4_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine4_syncfifo4_we;
wire hdmi2usbsoc_sdram_bankmachine4_syncfifo4_writable;
wire hdmi2usbsoc_sdram_bankmachine4_syncfifo4_re;
wire hdmi2usbsoc_sdram_bankmachine4_syncfifo4_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine4_syncfifo4_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine4_syncfifo4_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine4_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine4_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine4_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine4_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine4_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine4_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine4_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine4_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine4_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine4_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine4_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine4_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine4_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine4_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine4_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine4_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine4_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine4_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine4_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine4_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine4_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine4_hit;
reg hdmi2usbsoc_sdram_bankmachine4_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine4_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine4_wait;
wire hdmi2usbsoc_sdram_bankmachine4_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine4_count = 3'd4;
wire hdmi2usbsoc_sdram_bankmachine5_req_valid;
wire hdmi2usbsoc_sdram_bankmachine5_req_ready;
wire hdmi2usbsoc_sdram_bankmachine5_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine5_req_adr;
wire hdmi2usbsoc_sdram_bankmachine5_req_lock;
reg hdmi2usbsoc_sdram_bankmachine5_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine5_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine5_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine5_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine5_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine5_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine5_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine5_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine5_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine5_source_valid;
wire hdmi2usbsoc_sdram_bankmachine5_source_ready;
wire hdmi2usbsoc_sdram_bankmachine5_source_first;
wire hdmi2usbsoc_sdram_bankmachine5_source_last;
wire hdmi2usbsoc_sdram_bankmachine5_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine5_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine5_syncfifo5_we;
wire hdmi2usbsoc_sdram_bankmachine5_syncfifo5_writable;
wire hdmi2usbsoc_sdram_bankmachine5_syncfifo5_re;
wire hdmi2usbsoc_sdram_bankmachine5_syncfifo5_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine5_syncfifo5_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine5_syncfifo5_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine5_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine5_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine5_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine5_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine5_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine5_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine5_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine5_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine5_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine5_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine5_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine5_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine5_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine5_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine5_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine5_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine5_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine5_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine5_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine5_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine5_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine5_hit;
reg hdmi2usbsoc_sdram_bankmachine5_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine5_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine5_wait;
wire hdmi2usbsoc_sdram_bankmachine5_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine5_count = 3'd4;
wire hdmi2usbsoc_sdram_bankmachine6_req_valid;
wire hdmi2usbsoc_sdram_bankmachine6_req_ready;
wire hdmi2usbsoc_sdram_bankmachine6_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine6_req_adr;
wire hdmi2usbsoc_sdram_bankmachine6_req_lock;
reg hdmi2usbsoc_sdram_bankmachine6_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine6_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine6_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine6_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine6_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine6_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine6_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine6_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine6_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine6_source_valid;
wire hdmi2usbsoc_sdram_bankmachine6_source_ready;
wire hdmi2usbsoc_sdram_bankmachine6_source_first;
wire hdmi2usbsoc_sdram_bankmachine6_source_last;
wire hdmi2usbsoc_sdram_bankmachine6_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine6_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine6_syncfifo6_we;
wire hdmi2usbsoc_sdram_bankmachine6_syncfifo6_writable;
wire hdmi2usbsoc_sdram_bankmachine6_syncfifo6_re;
wire hdmi2usbsoc_sdram_bankmachine6_syncfifo6_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine6_syncfifo6_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine6_syncfifo6_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine6_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine6_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine6_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine6_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine6_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine6_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine6_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine6_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine6_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine6_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine6_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine6_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine6_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine6_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine6_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine6_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine6_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine6_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine6_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine6_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine6_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine6_hit;
reg hdmi2usbsoc_sdram_bankmachine6_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine6_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine6_wait;
wire hdmi2usbsoc_sdram_bankmachine6_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine6_count = 3'd4;
wire hdmi2usbsoc_sdram_bankmachine7_req_valid;
wire hdmi2usbsoc_sdram_bankmachine7_req_ready;
wire hdmi2usbsoc_sdram_bankmachine7_req_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine7_req_adr;
wire hdmi2usbsoc_sdram_bankmachine7_req_lock;
reg hdmi2usbsoc_sdram_bankmachine7_req_wdata_ready = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_req_rdata_valid = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine7_refresh_req;
reg hdmi2usbsoc_sdram_bankmachine7_refresh_gnt = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_ready = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine7_cmd_payload_a = 13'd0;
wire [2:0] hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ba;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_payload_we = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine7_sink_valid;
wire hdmi2usbsoc_sdram_bankmachine7_sink_ready;
reg hdmi2usbsoc_sdram_bankmachine7_sink_first = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_sink_last = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine7_sink_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine7_sink_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine7_source_valid;
wire hdmi2usbsoc_sdram_bankmachine7_source_ready;
wire hdmi2usbsoc_sdram_bankmachine7_source_first;
wire hdmi2usbsoc_sdram_bankmachine7_source_last;
wire hdmi2usbsoc_sdram_bankmachine7_source_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine7_source_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine7_syncfifo7_we;
wire hdmi2usbsoc_sdram_bankmachine7_syncfifo7_writable;
wire hdmi2usbsoc_sdram_bankmachine7_syncfifo7_re;
wire hdmi2usbsoc_sdram_bankmachine7_syncfifo7_readable;
wire [23:0] hdmi2usbsoc_sdram_bankmachine7_syncfifo7_din;
wire [23:0] hdmi2usbsoc_sdram_bankmachine7_syncfifo7_dout;
reg [3:0] hdmi2usbsoc_sdram_bankmachine7_level = 4'd0;
reg hdmi2usbsoc_sdram_bankmachine7_replace = 1'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine7_produce = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine7_consume = 3'd0;
reg [2:0] hdmi2usbsoc_sdram_bankmachine7_wrport_adr = 3'd0;
wire [23:0] hdmi2usbsoc_sdram_bankmachine7_wrport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine7_wrport_we;
wire [23:0] hdmi2usbsoc_sdram_bankmachine7_wrport_dat_w;
wire hdmi2usbsoc_sdram_bankmachine7_do_read;
wire [2:0] hdmi2usbsoc_sdram_bankmachine7_rdport_adr;
wire [23:0] hdmi2usbsoc_sdram_bankmachine7_rdport_dat_r;
wire hdmi2usbsoc_sdram_bankmachine7_fifo_in_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine7_fifo_in_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine7_fifo_in_first;
wire hdmi2usbsoc_sdram_bankmachine7_fifo_in_last;
wire hdmi2usbsoc_sdram_bankmachine7_fifo_out_payload_we;
wire [20:0] hdmi2usbsoc_sdram_bankmachine7_fifo_out_payload_adr;
wire hdmi2usbsoc_sdram_bankmachine7_fifo_out_first;
wire hdmi2usbsoc_sdram_bankmachine7_fifo_out_last;
reg hdmi2usbsoc_sdram_bankmachine7_has_openrow = 1'd0;
reg [12:0] hdmi2usbsoc_sdram_bankmachine7_openrow = 13'd0;
wire hdmi2usbsoc_sdram_bankmachine7_hit;
reg hdmi2usbsoc_sdram_bankmachine7_track_open = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_track_close = 1'd0;
reg hdmi2usbsoc_sdram_bankmachine7_sel_row_adr = 1'd0;
wire hdmi2usbsoc_sdram_bankmachine7_wait;
wire hdmi2usbsoc_sdram_bankmachine7_done;
reg [2:0] hdmi2usbsoc_sdram_bankmachine7_count = 3'd4;
reg hdmi2usbsoc_sdram_choose_cmd_want_reads = 1'd0;
reg hdmi2usbsoc_sdram_choose_cmd_want_writes = 1'd0;
reg hdmi2usbsoc_sdram_choose_cmd_want_cmds = 1'd0;
wire hdmi2usbsoc_sdram_choose_cmd_cmd_valid;
reg hdmi2usbsoc_sdram_choose_cmd_cmd_ready = 1'd0;
wire [12:0] hdmi2usbsoc_sdram_choose_cmd_cmd_payload_a;
wire [2:0] hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ba;
reg hdmi2usbsoc_sdram_choose_cmd_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_choose_cmd_cmd_payload_we = 1'd0;
wire hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_cmd;
wire hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_read;
wire hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_write;
reg [7:0] hdmi2usbsoc_sdram_choose_cmd_valids = 8'd0;
wire [7:0] hdmi2usbsoc_sdram_choose_cmd_request;
reg [2:0] hdmi2usbsoc_sdram_choose_cmd_grant = 3'd0;
wire hdmi2usbsoc_sdram_choose_cmd_ce;
reg hdmi2usbsoc_sdram_choose_req_want_reads = 1'd0;
reg hdmi2usbsoc_sdram_choose_req_want_writes = 1'd0;
reg hdmi2usbsoc_sdram_choose_req_want_cmds = 1'd0;
wire hdmi2usbsoc_sdram_choose_req_cmd_valid;
reg hdmi2usbsoc_sdram_choose_req_cmd_ready = 1'd0;
wire [12:0] hdmi2usbsoc_sdram_choose_req_cmd_payload_a;
wire [2:0] hdmi2usbsoc_sdram_choose_req_cmd_payload_ba;
reg hdmi2usbsoc_sdram_choose_req_cmd_payload_cas = 1'd0;
reg hdmi2usbsoc_sdram_choose_req_cmd_payload_ras = 1'd0;
reg hdmi2usbsoc_sdram_choose_req_cmd_payload_we = 1'd0;
wire hdmi2usbsoc_sdram_choose_req_cmd_payload_is_cmd;
wire hdmi2usbsoc_sdram_choose_req_cmd_payload_is_read;
wire hdmi2usbsoc_sdram_choose_req_cmd_payload_is_write;
reg [7:0] hdmi2usbsoc_sdram_choose_req_valids = 8'd0;
wire [7:0] hdmi2usbsoc_sdram_choose_req_request;
reg [2:0] hdmi2usbsoc_sdram_choose_req_grant = 3'd0;
wire hdmi2usbsoc_sdram_choose_req_ce;
reg [12:0] hdmi2usbsoc_sdram_nop_a = 13'd0;
reg [2:0] hdmi2usbsoc_sdram_nop_ba = 3'd0;
reg hdmi2usbsoc_sdram_nop_cas = 1'd0;
reg hdmi2usbsoc_sdram_nop_ras = 1'd0;
reg hdmi2usbsoc_sdram_nop_we = 1'd0;
reg [1:0] hdmi2usbsoc_sdram_sel0 = 2'd0;
reg [1:0] hdmi2usbsoc_sdram_sel1 = 2'd0;
wire hdmi2usbsoc_sdram_read_available;
wire hdmi2usbsoc_sdram_write_available;
reg hdmi2usbsoc_sdram_en0 = 1'd0;
wire hdmi2usbsoc_sdram_max_time0;
reg [4:0] hdmi2usbsoc_sdram_time0 = 5'd0;
reg hdmi2usbsoc_sdram_en1 = 1'd0;
wire hdmi2usbsoc_sdram_max_time1;
reg [3:0] hdmi2usbsoc_sdram_time1 = 4'd0;
wire hdmi2usbsoc_sdram_go_to_refresh;
wire hdmi2usbsoc_sdram_bandwidth_update_re;
wire hdmi2usbsoc_sdram_bandwidth_update_r;
reg hdmi2usbsoc_sdram_bandwidth_update_w = 1'd0;
reg [23:0] hdmi2usbsoc_sdram_bandwidth_nreads_status = 24'd0;
reg [23:0] hdmi2usbsoc_sdram_bandwidth_nwrites_status = 24'd0;
reg [6:0] hdmi2usbsoc_sdram_bandwidth_data_width_status = 7'd64;
reg hdmi2usbsoc_sdram_bandwidth_cmd_valid = 1'd0;
reg hdmi2usbsoc_sdram_bandwidth_cmd_ready = 1'd0;
reg hdmi2usbsoc_sdram_bandwidth_cmd_is_read = 1'd0;
reg hdmi2usbsoc_sdram_bandwidth_cmd_is_write = 1'd0;
reg [23:0] hdmi2usbsoc_sdram_bandwidth_counter = 24'd0;
reg hdmi2usbsoc_sdram_bandwidth_period = 1'd0;
reg [23:0] hdmi2usbsoc_sdram_bandwidth_nreads = 24'd0;
reg [23:0] hdmi2usbsoc_sdram_bandwidth_nwrites = 24'd0;
reg [23:0] hdmi2usbsoc_sdram_bandwidth_nreads_r = 24'd0;
reg [23:0] hdmi2usbsoc_sdram_bandwidth_nwrites_r = 24'd0;
wire [29:0] hdmi2usbsoc_interface1_wb_sdram_adr;
wire [31:0] hdmi2usbsoc_interface1_wb_sdram_dat_w;
wire [31:0] hdmi2usbsoc_interface1_wb_sdram_dat_r;
wire [3:0] hdmi2usbsoc_interface1_wb_sdram_sel;
wire hdmi2usbsoc_interface1_wb_sdram_cyc;
wire hdmi2usbsoc_interface1_wb_sdram_stb;
wire hdmi2usbsoc_interface1_wb_sdram_ack;
wire hdmi2usbsoc_interface1_wb_sdram_we;
wire [2:0] hdmi2usbsoc_interface1_wb_sdram_cti;
wire [1:0] hdmi2usbsoc_interface1_wb_sdram_bte;
wire hdmi2usbsoc_interface1_wb_sdram_err;
reg hdmi2usbsoc_port_cmd_valid = 1'd0;
wire hdmi2usbsoc_port_cmd_ready;
reg hdmi2usbsoc_port_cmd_payload_we = 1'd0;
wire [23:0] hdmi2usbsoc_port_cmd_payload_adr;
reg hdmi2usbsoc_port_wdata_valid = 1'd0;
wire hdmi2usbsoc_port_wdata_ready;
wire [63:0] hdmi2usbsoc_port_wdata_payload_data;
wire [7:0] hdmi2usbsoc_port_wdata_payload_we;
wire hdmi2usbsoc_port_rdata_valid;
reg hdmi2usbsoc_port_rdata_ready = 1'd0;
wire [63:0] hdmi2usbsoc_port_rdata_payload_data;
wire [29:0] hdmi2usbsoc_interface_adr;
wire [63:0] hdmi2usbsoc_interface_dat_w;
wire [63:0] hdmi2usbsoc_interface_dat_r;
wire [7:0] hdmi2usbsoc_interface_sel;
reg hdmi2usbsoc_interface_cyc = 1'd0;
reg hdmi2usbsoc_interface_stb = 1'd0;
reg hdmi2usbsoc_interface_ack = 1'd0;
reg hdmi2usbsoc_interface_we = 1'd0;
wire [9:0] hdmi2usbsoc_data_port_adr;
wire [63:0] hdmi2usbsoc_data_port_dat_r;
reg [7:0] hdmi2usbsoc_data_port_we = 8'd0;
reg [63:0] hdmi2usbsoc_data_port_dat_w = 64'd0;
reg hdmi2usbsoc_write_from_slave = 1'd0;
reg hdmi2usbsoc_adr_offset_r = 1'd0;
wire [9:0] hdmi2usbsoc_tag_port_adr;
wire [21:0] hdmi2usbsoc_tag_port_dat_r;
reg hdmi2usbsoc_tag_port_we = 1'd0;
wire [21:0] hdmi2usbsoc_tag_port_dat_w;
wire [20:0] hdmi2usbsoc_tag_do_tag;
wire hdmi2usbsoc_tag_do_dirty;
wire [20:0] hdmi2usbsoc_tag_di_tag;
reg hdmi2usbsoc_tag_di_dirty = 1'd0;
reg hdmi2usbsoc_word_clr = 1'd0;
reg hdmi2usbsoc_word_inc = 1'd0;
wire hdmi2usbsoc_litedramport0_cmd_valid0;
wire hdmi2usbsoc_litedramport0_cmd_ready0;
wire hdmi2usbsoc_litedramport0_cmd_payload_we0;
wire [23:0] hdmi2usbsoc_litedramport0_cmd_payload_adr0;
wire hdmi2usbsoc_litedramport0_wdata_valid;
wire hdmi2usbsoc_litedramport0_wdata_ready;
wire [63:0] hdmi2usbsoc_litedramport0_wdata_payload_data;
wire [7:0] hdmi2usbsoc_litedramport0_wdata_payload_we;
wire hdmi2usbsoc_litedramport0_rdata_valid0;
wire [63:0] hdmi2usbsoc_litedramport0_rdata_payload_data0;
wire hdmi2usbsoc_hdmi_in0_edid_status;
reg hdmi2usbsoc_hdmi_in0_edid_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi_in0_edid_storage;
reg hdmi2usbsoc_hdmi_in0_edid_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_edid_scl_raw;
reg hdmi2usbsoc_hdmi_in0_edid_sda_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_edid_sda_raw;
reg hdmi2usbsoc_hdmi_in0_edid_sda_drv = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_sda_drv_reg = 1'd0;
wire hdmi2usbsoc_hdmi_in0_edid_sda_i_async;
wire hdmi2usbsoc_hdmi_in0_edid_sda_o;
reg hdmi2usbsoc_hdmi_in0_edid_scl_i = 1'd0;
reg [5:0] hdmi2usbsoc_hdmi_in0_edid_samp_count = 6'd0;
reg hdmi2usbsoc_hdmi_in0_edid_samp_carry = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_scl_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_sda_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_edid_scl_rising;
wire hdmi2usbsoc_hdmi_in0_edid_sda_rising;
wire hdmi2usbsoc_hdmi_in0_edid_sda_falling;
wire hdmi2usbsoc_hdmi_in0_edid_start;
reg [7:0] hdmi2usbsoc_hdmi_in0_edid_din = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_edid_counter = 4'd0;
reg hdmi2usbsoc_hdmi_in0_edid_is_read = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_update_is_read = 1'd0;
reg [6:0] hdmi2usbsoc_hdmi_in0_edid_offset_counter = 7'd0;
reg hdmi2usbsoc_hdmi_in0_edid_oc_load = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_oc_inc = 1'd0;
wire [6:0] hdmi2usbsoc_hdmi_in0_edid_adr;
wire [7:0] hdmi2usbsoc_hdmi_in0_edid_dat_r;
reg hdmi2usbsoc_hdmi_in0_edid_data_bit = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_zero_drv = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_data_drv = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_data_drv_en = 1'd0;
reg hdmi2usbsoc_hdmi_in0_edid_data_drv_stop = 1'd0;
reg hdmi2usbsoc_hdmi_in0_pll_reset_storage_full = 1'd1;
wire hdmi2usbsoc_hdmi_in0_pll_reset_storage;
reg hdmi2usbsoc_hdmi_in0_pll_reset_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_locked_status;
reg [4:0] hdmi2usbsoc_hdmi_in0_pll_adr_storage_full = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_in0_pll_adr_storage;
reg hdmi2usbsoc_hdmi_in0_pll_adr_re = 1'd0;
wire [15:0] hdmi2usbsoc_hdmi_in0_pll_dat_r_status;
reg [15:0] hdmi2usbsoc_hdmi_in0_pll_dat_w_storage_full = 16'd0;
wire [15:0] hdmi2usbsoc_hdmi_in0_pll_dat_w_storage;
reg hdmi2usbsoc_hdmi_in0_pll_dat_w_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_pll_read_re;
wire hdmi2usbsoc_hdmi_in0_pll_read_r;
reg hdmi2usbsoc_hdmi_in0_pll_read_w = 1'd0;
wire hdmi2usbsoc_hdmi_in0_pll_write_re;
wire hdmi2usbsoc_hdmi_in0_pll_write_r;
reg hdmi2usbsoc_hdmi_in0_pll_write_w = 1'd0;
reg hdmi2usbsoc_hdmi_in0_pll_drdy_status = 1'd0;
wire hdmi2usbsoc_hdmi_in0_locked;
wire hdmi2usbsoc_hdmi_in0_serdesstrobe;
wire hdmi_in0_pix_clk;
wire hdmi_in0_pix_rst;
wire hdmi_in0_pix_o_clk;
reg hdmi_in0_pix_o_rst = 1'd0;
wire hdmi_in0_pix2x_clk;
wire hdmi_in0_pix2x_rst;
wire hdmi_in0_pix10x_clk;
wire hdmi2usbsoc_hdmi_in0_clk_input;
wire hdmi2usbsoc_hdmi_in0_clkfbout;
wire hdmi2usbsoc_hdmi_in0_pll_locked;
wire hdmi2usbsoc_hdmi_in0_pll_clk0;
wire hdmi2usbsoc_hdmi_in0_pll_clk1;
wire hdmi2usbsoc_hdmi_in0_pll_clk2;
wire hdmi2usbsoc_hdmi_in0_pll_drdy;
wire hdmi2usbsoc_hdmi_in0_locked_async;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_serdesstrobe;
reg [9:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_d = 10'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re;
wire [5:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r;
reg [5:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_w = 6'd0;
wire [1:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_busy_status;
wire [1:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_status;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_reset_re;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_reset_r;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_reset_w = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_se;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_delayed_master;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_delayed_slave;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_inc;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_ce;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_cal;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_rst;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_busy;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_cal;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_rst;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_busy;
wire [4:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr2;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_valid;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_incdec;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_edge;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_cascade;
reg [7:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness = 8'd128;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_too_late;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_too_early;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_reset_lateness;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_o_r = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_charsync0_raw_data;
reg hdmi2usbsoc_hdmi_in0_charsync0_synced = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_charsync0_data = 10'd0;
wire hdmi2usbsoc_hdmi_in0_charsync0_char_synced_status;
wire [3:0] hdmi2usbsoc_hdmi_in0_charsync0_ctl_pos_status;
reg [9:0] hdmi2usbsoc_hdmi_in0_charsync0_raw_data1 = 10'd0;
wire [19:0] hdmi2usbsoc_hdmi_in0_charsync0_raw;
reg hdmi2usbsoc_hdmi_in0_charsync0_found_control = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync0_control_position = 4'd0;
reg [2:0] hdmi2usbsoc_hdmi_in0_charsync0_control_counter = 3'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync0_previous_control_position = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync0_word_sel = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_wer0_data;
wire hdmi2usbsoc_hdmi_in0_wer0_update_re;
wire hdmi2usbsoc_hdmi_in0_wer0_update_r;
reg hdmi2usbsoc_hdmi_in0_wer0_update_w = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer0_status = 24'd0;
reg [8:0] hdmi2usbsoc_hdmi_in0_wer0_data_r = 9'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_wer0_transitions = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_wer0_transition_count = 4'd0;
reg hdmi2usbsoc_hdmi_in0_wer0_is_control = 1'd0;
reg hdmi2usbsoc_hdmi_in0_wer0_is_error = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer0_period_counter = 24'd0;
reg hdmi2usbsoc_hdmi_in0_wer0_period_done = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer0_wer_counter = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r = 24'd0;
reg hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r_updated = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer0_wer_counter_sys = 24'd0;
wire hdmi2usbsoc_hdmi_in0_wer0_i;
wire hdmi2usbsoc_hdmi_in0_wer0_o;
reg hdmi2usbsoc_hdmi_in0_wer0_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_wer0_toggle_o;
reg hdmi2usbsoc_hdmi_in0_wer0_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_decoding0_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in0_decoding0_input;
reg hdmi2usbsoc_hdmi_in0_decoding0_valid_o = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_decoding0_output_raw = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_decoding0_output_d = 8'd0;
reg [1:0] hdmi2usbsoc_hdmi_in0_decoding0_output_c = 2'd0;
reg hdmi2usbsoc_hdmi_in0_decoding0_output_de = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_serdesstrobe;
reg [9:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_d = 10'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re;
wire [5:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r;
reg [5:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_w = 6'd0;
wire [1:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_busy_status;
wire [1:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_status;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_reset_re;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_reset_r;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_reset_w = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_se;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_delayed_master;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_delayed_slave;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_inc;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_ce;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_cal;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_rst;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_busy;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_cal;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_rst;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_busy;
wire [4:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr2;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_valid;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_incdec;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_edge;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_cascade;
reg [7:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness = 8'd128;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_too_late;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_too_early;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_reset_lateness;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_o_r = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_charsync1_raw_data;
reg hdmi2usbsoc_hdmi_in0_charsync1_synced = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_charsync1_data = 10'd0;
wire hdmi2usbsoc_hdmi_in0_charsync1_char_synced_status;
wire [3:0] hdmi2usbsoc_hdmi_in0_charsync1_ctl_pos_status;
reg [9:0] hdmi2usbsoc_hdmi_in0_charsync1_raw_data1 = 10'd0;
wire [19:0] hdmi2usbsoc_hdmi_in0_charsync1_raw;
reg hdmi2usbsoc_hdmi_in0_charsync1_found_control = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync1_control_position = 4'd0;
reg [2:0] hdmi2usbsoc_hdmi_in0_charsync1_control_counter = 3'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync1_previous_control_position = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync1_word_sel = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_wer1_data;
wire hdmi2usbsoc_hdmi_in0_wer1_update_re;
wire hdmi2usbsoc_hdmi_in0_wer1_update_r;
reg hdmi2usbsoc_hdmi_in0_wer1_update_w = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer1_status = 24'd0;
reg [8:0] hdmi2usbsoc_hdmi_in0_wer1_data_r = 9'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_wer1_transitions = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_wer1_transition_count = 4'd0;
reg hdmi2usbsoc_hdmi_in0_wer1_is_control = 1'd0;
reg hdmi2usbsoc_hdmi_in0_wer1_is_error = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer1_period_counter = 24'd0;
reg hdmi2usbsoc_hdmi_in0_wer1_period_done = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer1_wer_counter = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r = 24'd0;
reg hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r_updated = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer1_wer_counter_sys = 24'd0;
wire hdmi2usbsoc_hdmi_in0_wer1_i;
wire hdmi2usbsoc_hdmi_in0_wer1_o;
reg hdmi2usbsoc_hdmi_in0_wer1_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_wer1_toggle_o;
reg hdmi2usbsoc_hdmi_in0_wer1_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_decoding1_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in0_decoding1_input;
reg hdmi2usbsoc_hdmi_in0_decoding1_valid_o = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_decoding1_output_raw = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_decoding1_output_d = 8'd0;
reg [1:0] hdmi2usbsoc_hdmi_in0_decoding1_output_c = 2'd0;
reg hdmi2usbsoc_hdmi_in0_decoding1_output_de = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_serdesstrobe;
reg [9:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_d = 10'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re;
wire [5:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r;
reg [5:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_w = 6'd0;
wire [1:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_busy_status;
wire [1:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_status;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_reset_re;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_reset_r;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_reset_w = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_se;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_delayed_master;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_delayed_slave;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_inc;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_ce;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_cal;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_rst;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_busy;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_cal;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_rst;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_busy;
wire [4:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr2;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_valid;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_incdec;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_edge;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_cascade;
reg [7:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness = 8'd128;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_too_late;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_too_early;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_reset_lateness;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_i;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_o;
reg hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_o_r = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_charsync2_raw_data;
reg hdmi2usbsoc_hdmi_in0_charsync2_synced = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_charsync2_data = 10'd0;
wire hdmi2usbsoc_hdmi_in0_charsync2_char_synced_status;
wire [3:0] hdmi2usbsoc_hdmi_in0_charsync2_ctl_pos_status;
reg [9:0] hdmi2usbsoc_hdmi_in0_charsync2_raw_data1 = 10'd0;
wire [19:0] hdmi2usbsoc_hdmi_in0_charsync2_raw;
reg hdmi2usbsoc_hdmi_in0_charsync2_found_control = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync2_control_position = 4'd0;
reg [2:0] hdmi2usbsoc_hdmi_in0_charsync2_control_counter = 3'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync2_previous_control_position = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_charsync2_word_sel = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_wer2_data;
wire hdmi2usbsoc_hdmi_in0_wer2_update_re;
wire hdmi2usbsoc_hdmi_in0_wer2_update_r;
reg hdmi2usbsoc_hdmi_in0_wer2_update_w = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer2_status = 24'd0;
reg [8:0] hdmi2usbsoc_hdmi_in0_wer2_data_r = 9'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_wer2_transitions = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_wer2_transition_count = 4'd0;
reg hdmi2usbsoc_hdmi_in0_wer2_is_control = 1'd0;
reg hdmi2usbsoc_hdmi_in0_wer2_is_error = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer2_period_counter = 24'd0;
reg hdmi2usbsoc_hdmi_in0_wer2_period_done = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer2_wer_counter = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r = 24'd0;
reg hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r_updated = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_wer2_wer_counter_sys = 24'd0;
wire hdmi2usbsoc_hdmi_in0_wer2_i;
wire hdmi2usbsoc_hdmi_in0_wer2_o;
reg hdmi2usbsoc_hdmi_in0_wer2_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_wer2_toggle_o;
reg hdmi2usbsoc_hdmi_in0_wer2_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_decoding2_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in0_decoding2_input;
reg hdmi2usbsoc_hdmi_in0_decoding2_valid_o = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_decoding2_output_raw = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_decoding2_output_d = 8'd0;
reg [1:0] hdmi2usbsoc_hdmi_in0_decoding2_output_c = 2'd0;
reg hdmi2usbsoc_hdmi_in0_decoding2_output_de = 1'd0;
wire hdmi2usbsoc_hdmi_in0_chansync_valid_i;
reg hdmi2usbsoc_hdmi_in0_chansync_chan_synced = 1'd0;
wire hdmi2usbsoc_hdmi_in0_chansync_status;
wire hdmi2usbsoc_hdmi_in0_chansync_all_control;
wire [9:0] hdmi2usbsoc_hdmi_in0_chansync_data_in0_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_chansync_data_in0_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_chansync_data_in0_c;
wire hdmi2usbsoc_hdmi_in0_chansync_data_in0_de;
wire [9:0] hdmi2usbsoc_hdmi_in0_chansync_data_out0_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_chansync_data_out0_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_chansync_data_out0_c;
wire hdmi2usbsoc_hdmi_in0_chansync_data_out0_de;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_din;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_dout;
wire hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_re;
reg [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_produce = 3'd0;
reg [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_consume = 3'd0;
wire [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_we;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_w;
wire [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_rdport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in0_chansync_is_control0;
wire [9:0] hdmi2usbsoc_hdmi_in0_chansync_data_in1_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_chansync_data_in1_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_chansync_data_in1_c;
wire hdmi2usbsoc_hdmi_in0_chansync_data_in1_de;
wire [9:0] hdmi2usbsoc_hdmi_in0_chansync_data_out1_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_chansync_data_out1_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_chansync_data_out1_c;
wire hdmi2usbsoc_hdmi_in0_chansync_data_out1_de;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_din;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_dout;
wire hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_re;
reg [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_produce = 3'd0;
reg [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_consume = 3'd0;
wire [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_we;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_w;
wire [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_rdport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in0_chansync_is_control1;
wire [9:0] hdmi2usbsoc_hdmi_in0_chansync_data_in2_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_chansync_data_in2_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_chansync_data_in2_c;
wire hdmi2usbsoc_hdmi_in0_chansync_data_in2_de;
wire [9:0] hdmi2usbsoc_hdmi_in0_chansync_data_out2_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_chansync_data_out2_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_chansync_data_out2_c;
wire hdmi2usbsoc_hdmi_in0_chansync_data_out2_de;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_din;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_dout;
wire hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_re;
reg [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_produce = 3'd0;
reg [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_consume = 3'd0;
wire [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_we;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_w;
wire [2:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_rdport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in0_chansync_is_control2;
wire hdmi2usbsoc_hdmi_in0_chansync_some_control;
wire hdmi2usbsoc_hdmi_in0_syncpol_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in0_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in0_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in0_c;
wire hdmi2usbsoc_hdmi_in0_syncpol_data_in0_de;
wire [9:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in1_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in1_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in1_c;
wire hdmi2usbsoc_hdmi_in0_syncpol_data_in1_de;
wire [9:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in2_raw;
wire [7:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in2_d;
wire [1:0] hdmi2usbsoc_hdmi_in0_syncpol_data_in2_c;
wire hdmi2usbsoc_hdmi_in0_syncpol_data_in2_de;
reg hdmi2usbsoc_hdmi_in0_syncpol_valid_o = 1'd0;
wire hdmi2usbsoc_hdmi_in0_syncpol_de;
wire hdmi2usbsoc_hdmi_in0_syncpol_hsync;
wire hdmi2usbsoc_hdmi_in0_syncpol_vsync;
reg [7:0] hdmi2usbsoc_hdmi_in0_syncpol_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_syncpol_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_syncpol_b = 8'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_syncpol_c0 = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_syncpol_c1 = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_syncpol_c2 = 10'd0;
reg hdmi2usbsoc_hdmi_in0_syncpol_de_r = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_in0_syncpol_c_polarity = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_in0_syncpol_c_out = 2'd0;
wire hdmi2usbsoc_hdmi_in0_resdetection_valid_i;
wire hdmi2usbsoc_hdmi_in0_resdetection_vsync;
wire hdmi2usbsoc_hdmi_in0_resdetection_de;
wire [10:0] hdmi2usbsoc_hdmi_in0_resdetection_hres_status;
wire [10:0] hdmi2usbsoc_hdmi_in0_resdetection_vres_status;
reg hdmi2usbsoc_hdmi_in0_resdetection_de_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_resdetection_pn_de;
reg [10:0] hdmi2usbsoc_hdmi_in0_resdetection_hcounter = 11'd0;
reg [10:0] hdmi2usbsoc_hdmi_in0_resdetection_hcounter_st = 11'd0;
reg hdmi2usbsoc_hdmi_in0_resdetection_vsync_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_resdetection_p_vsync;
reg [10:0] hdmi2usbsoc_hdmi_in0_resdetection_vcounter = 11'd0;
reg [10:0] hdmi2usbsoc_hdmi_in0_resdetection_vcounter_st = 11'd0;
wire hdmi2usbsoc_hdmi_in0_frame_valid_i;
wire hdmi2usbsoc_hdmi_in0_frame_vsync;
wire hdmi2usbsoc_hdmi_in0_frame_de;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_r;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_g;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_b;
wire hdmi2usbsoc_hdmi_in0_frame_frame_valid;
wire hdmi2usbsoc_hdmi_in0_frame_frame_ready;
wire hdmi2usbsoc_hdmi_in0_frame_frame_first;
wire hdmi2usbsoc_hdmi_in0_frame_frame_last;
wire hdmi2usbsoc_hdmi_in0_frame_frame_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in0_frame_frame_payload_pixels;
wire hdmi2usbsoc_hdmi_in0_frame_busy;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_re;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_r;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_w;
reg hdmi2usbsoc_hdmi_in0_frame_de_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_valid;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_ready;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_last = 1'd0;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_b;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_valid;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_ready;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_first;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_last;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_cr;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_r;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_g;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_b;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_b = 8'd0;
reg signed [8:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_g = 9'sd0;
reg signed [8:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_g = 9'sd0;
reg signed [16:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_ca_mult_rg = 17'sd0;
reg signed [16:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb_mult_bg = 17'sd0;
reg signed [24:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_carg_plus_cbbg = 25'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw = 11'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_yraw = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_yraw = 12'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r0 = 11'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cc_mult_ryraw = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cd_mult_byraw = 20'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r1 = 11'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_y = 11'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cr = 12'sd0;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_ce;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce;
wire hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_busy;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n4 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n5 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n6 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n7 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n4 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n4 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n5 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n5 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n6 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n6 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n7 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n7 = 1'd0;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_valid;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_ready;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_first;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_cr;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_valid;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_ready;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_first;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_last;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_payload_cb_cr;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_y;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cb;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cr;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_cb_cr = 8'd0;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_cr = 8'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_parity = 1'd0;
reg [8:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cb_sum = 9'd0;
reg [8:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cr_sum = 9'd0;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cb_mean;
wire [7:0] hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cr_mean;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_ce;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce;
wire hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_busy;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync0 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync1 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync2 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de3 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync3 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de4 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync4 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de5 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync5 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de6 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync6 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de7 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync7 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de8 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync8 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de9 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync9 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_de10 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_next_vsync10 = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_vsync_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_frame_new_frame;
reg [63:0] hdmi2usbsoc_hdmi_in0_frame_cur_word = 64'd0;
reg hdmi2usbsoc_hdmi_in0_frame_cur_word_valid = 1'd0;
wire [15:0] hdmi2usbsoc_hdmi_in0_frame_encoded_pixel;
reg [1:0] hdmi2usbsoc_hdmi_in0_frame_pack_counter = 2'd0;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_sink_valid;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_in0_frame_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_fifo_sink_last = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_sof = 1'd0;
wire [63:0] hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_pixels;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_source_valid;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_source_ready;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_source_first;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_source_last;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_source_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in0_frame_fifo_source_payload_pixels;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_we;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_writable;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_re;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_readable;
wire [66:0] hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_din;
wire [66:0] hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_dout;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_ce;
(* register_balancing = "no" *) reg [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next;
reg [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_binary = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next_binary = 10'd0;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_ce;
(* register_balancing = "no" *) reg [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next;
reg [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_binary = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_produce_rdomain;
wire [9:0] hdmi2usbsoc_hdmi_in0_frame_fifo_consume_wdomain;
wire [8:0] hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_adr;
wire [66:0] hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_we;
wire [66:0] hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_dat_w;
wire [8:0] hdmi2usbsoc_hdmi_in0_frame_fifo_rdport_adr;
wire [66:0] hdmi2usbsoc_hdmi_in0_frame_fifo_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_payload_pixels;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_last;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_payload_pixels;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_in0_frame_pix_overflow = 1'd0;
wire hdmi2usbsoc_hdmi_in0_frame_pix_overflow_reset;
wire hdmi2usbsoc_hdmi_in0_frame_sys_overflow;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_reset_i;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_reset_o;
reg hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_o;
reg hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_i;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_o;
reg hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_o;
reg hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in0_frame_overflow_mask = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_frame_valid;
reg hdmi2usbsoc_hdmi_in0_dma_frame_ready = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_frame_first;
wire hdmi2usbsoc_hdmi_in0_dma_frame_last;
wire hdmi2usbsoc_hdmi_in0_dma_frame_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in0_dma_frame_payload_pixels;
reg [26:0] hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full = 27'd0;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_frame_size_storage;
reg hdmi2usbsoc_hdmi_in0_dma_frame_size_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_irq;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_address;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_address_reached;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_address_valid;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_address_done = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_pending;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_trigger;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_clear = 1'd0;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_reached;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_valid;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_done;
reg [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage_full = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_we;
wire [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_dat_w;
reg [26:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full = 27'd0;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_we;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_dat_w;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_pending;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_trigger;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_clear = 1'd0;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_reached;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_valid;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_done;
reg [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage_full = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_we;
wire [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_dat_w;
reg [26:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full = 27'd0;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_we;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_dat_w;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_status_re;
wire [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_status_r;
reg [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_status_w = 2'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_re;
wire [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_r;
reg [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_w = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_storage_full = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_in0_dma_slot_array_storage;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_re = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_slot_array_change_slot;
reg hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot = 1'd0;
reg hdmi2usbsoc_hdmi_in0_dma_reset_words = 1'd0;
reg hdmi2usbsoc_hdmi_in0_dma_count_word = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_last_word;
reg [23:0] hdmi2usbsoc_hdmi_in0_dma_current_address = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in0_dma_mwords_remaining = 24'd0;
wire [63:0] hdmi2usbsoc_hdmi_in0_dma_memory_word;
reg hdmi2usbsoc_hdmi_in0_dma_sink_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_in0_dma_sink_sink_ready;
wire [23:0] hdmi2usbsoc_hdmi_in0_dma_sink_sink_payload_address;
wire [63:0] hdmi2usbsoc_hdmi_in0_dma_sink_sink_payload_data;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_sink_valid;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_in0_dma_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_in0_dma_fifo_sink_last = 1'd0;
wire [63:0] hdmi2usbsoc_hdmi_in0_dma_fifo_sink_payload_data;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_source_valid;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_source_ready;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_source_first;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_source_last;
wire [63:0] hdmi2usbsoc_hdmi_in0_dma_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_readable;
wire [65:0] hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_din;
wire [65:0] hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_dout;
reg [4:0] hdmi2usbsoc_hdmi_in0_dma_fifo_level = 5'd0;
reg hdmi2usbsoc_hdmi_in0_dma_fifo_replace = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_dma_fifo_produce = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_dma_fifo_consume = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_adr = 4'd0;
wire [65:0] hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_we;
wire [65:0] hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_do_read;
wire [3:0] hdmi2usbsoc_hdmi_in0_dma_fifo_rdport_adr;
wire [65:0] hdmi2usbsoc_hdmi_in0_dma_fifo_rdport_dat_r;
wire [63:0] hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_last;
wire [63:0] hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_last;
wire hdmi2usbsoc_litedramport1_cmd_valid0;
wire hdmi2usbsoc_litedramport1_cmd_ready0;
wire hdmi2usbsoc_litedramport1_cmd_payload_we0;
wire [23:0] hdmi2usbsoc_litedramport1_cmd_payload_adr0;
wire hdmi2usbsoc_litedramport1_wdata_valid;
wire hdmi2usbsoc_litedramport1_wdata_ready;
wire [63:0] hdmi2usbsoc_litedramport1_wdata_payload_data;
wire [7:0] hdmi2usbsoc_litedramport1_wdata_payload_we;
wire hdmi2usbsoc_litedramport1_rdata_valid0;
wire [63:0] hdmi2usbsoc_litedramport1_rdata_payload_data0;
wire hdmi2usbsoc_hdmi_in1_edid_status;
reg hdmi2usbsoc_hdmi_in1_edid_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi_in1_edid_storage;
reg hdmi2usbsoc_hdmi_in1_edid_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_edid_scl_raw;
reg hdmi2usbsoc_hdmi_in1_edid_sda_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_edid_sda_raw;
reg hdmi2usbsoc_hdmi_in1_edid_sda_drv = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_sda_drv_reg = 1'd0;
wire hdmi2usbsoc_hdmi_in1_edid_sda_i_async;
wire hdmi2usbsoc_hdmi_in1_edid_sda_o;
reg hdmi2usbsoc_hdmi_in1_edid_scl_i = 1'd0;
reg [5:0] hdmi2usbsoc_hdmi_in1_edid_samp_count = 6'd0;
reg hdmi2usbsoc_hdmi_in1_edid_samp_carry = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_scl_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_sda_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_edid_scl_rising;
wire hdmi2usbsoc_hdmi_in1_edid_sda_rising;
wire hdmi2usbsoc_hdmi_in1_edid_sda_falling;
wire hdmi2usbsoc_hdmi_in1_edid_start;
reg [7:0] hdmi2usbsoc_hdmi_in1_edid_din = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_edid_counter = 4'd0;
reg hdmi2usbsoc_hdmi_in1_edid_is_read = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_update_is_read = 1'd0;
reg [6:0] hdmi2usbsoc_hdmi_in1_edid_offset_counter = 7'd0;
reg hdmi2usbsoc_hdmi_in1_edid_oc_load = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_oc_inc = 1'd0;
wire [6:0] hdmi2usbsoc_hdmi_in1_edid_adr;
wire [7:0] hdmi2usbsoc_hdmi_in1_edid_dat_r;
reg hdmi2usbsoc_hdmi_in1_edid_data_bit = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_zero_drv = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_data_drv = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_data_drv_en = 1'd0;
reg hdmi2usbsoc_hdmi_in1_edid_data_drv_stop = 1'd0;
reg hdmi2usbsoc_hdmi_in1_pll_reset_storage_full = 1'd1;
wire hdmi2usbsoc_hdmi_in1_pll_reset_storage;
reg hdmi2usbsoc_hdmi_in1_pll_reset_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_locked_status;
reg [4:0] hdmi2usbsoc_hdmi_in1_pll_adr_storage_full = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_in1_pll_adr_storage;
reg hdmi2usbsoc_hdmi_in1_pll_adr_re = 1'd0;
wire [15:0] hdmi2usbsoc_hdmi_in1_pll_dat_r_status;
reg [15:0] hdmi2usbsoc_hdmi_in1_pll_dat_w_storage_full = 16'd0;
wire [15:0] hdmi2usbsoc_hdmi_in1_pll_dat_w_storage;
reg hdmi2usbsoc_hdmi_in1_pll_dat_w_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_pll_read_re;
wire hdmi2usbsoc_hdmi_in1_pll_read_r;
reg hdmi2usbsoc_hdmi_in1_pll_read_w = 1'd0;
wire hdmi2usbsoc_hdmi_in1_pll_write_re;
wire hdmi2usbsoc_hdmi_in1_pll_write_r;
reg hdmi2usbsoc_hdmi_in1_pll_write_w = 1'd0;
reg hdmi2usbsoc_hdmi_in1_pll_drdy_status = 1'd0;
wire hdmi2usbsoc_hdmi_in1_locked;
wire hdmi2usbsoc_hdmi_in1_serdesstrobe;
wire hdmi_in1_pix_clk;
wire hdmi_in1_pix_rst;
wire hdmi_in1_pix_o_clk;
reg hdmi_in1_pix_o_rst = 1'd0;
wire hdmi_in1_pix2x_clk;
wire hdmi_in1_pix2x_rst;
wire hdmi_in1_pix10x_clk;
wire hdmi2usbsoc_hdmi_in1_clk_input;
wire hdmi2usbsoc_hdmi_in1_clkfbout;
wire hdmi2usbsoc_hdmi_in1_pll_locked;
wire hdmi2usbsoc_hdmi_in1_pll_clk0;
wire hdmi2usbsoc_hdmi_in1_pll_clk1;
wire hdmi2usbsoc_hdmi_in1_pll_clk2;
wire hdmi2usbsoc_hdmi_in1_pll_drdy;
wire hdmi2usbsoc_hdmi_in1_locked_async;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_serdesstrobe;
reg [9:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_d = 10'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re;
wire [5:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r;
reg [5:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_w = 6'd0;
wire [1:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_busy_status;
wire [1:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_status;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_reset_re;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_reset_r;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_reset_w = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_se;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_delayed_master;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_delayed_slave;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_inc;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_ce;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_cal;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_rst;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_busy;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_cal;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_rst;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_busy;
wire [4:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr2;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_valid;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_incdec;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_edge;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_cascade;
reg [7:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness = 8'd128;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_too_late;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_too_early;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_reset_lateness;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_o_r = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_charsync0_raw_data;
reg hdmi2usbsoc_hdmi_in1_charsync0_synced = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_charsync0_data = 10'd0;
wire hdmi2usbsoc_hdmi_in1_charsync0_char_synced_status;
wire [3:0] hdmi2usbsoc_hdmi_in1_charsync0_ctl_pos_status;
reg [9:0] hdmi2usbsoc_hdmi_in1_charsync0_raw_data1 = 10'd0;
wire [19:0] hdmi2usbsoc_hdmi_in1_charsync0_raw;
reg hdmi2usbsoc_hdmi_in1_charsync0_found_control = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync0_control_position = 4'd0;
reg [2:0] hdmi2usbsoc_hdmi_in1_charsync0_control_counter = 3'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync0_previous_control_position = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync0_word_sel = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_wer0_data;
wire hdmi2usbsoc_hdmi_in1_wer0_update_re;
wire hdmi2usbsoc_hdmi_in1_wer0_update_r;
reg hdmi2usbsoc_hdmi_in1_wer0_update_w = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer0_status = 24'd0;
reg [8:0] hdmi2usbsoc_hdmi_in1_wer0_data_r = 9'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_wer0_transitions = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_wer0_transition_count = 4'd0;
reg hdmi2usbsoc_hdmi_in1_wer0_is_control = 1'd0;
reg hdmi2usbsoc_hdmi_in1_wer0_is_error = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer0_period_counter = 24'd0;
reg hdmi2usbsoc_hdmi_in1_wer0_period_done = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer0_wer_counter = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r = 24'd0;
reg hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r_updated = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer0_wer_counter_sys = 24'd0;
wire hdmi2usbsoc_hdmi_in1_wer0_i;
wire hdmi2usbsoc_hdmi_in1_wer0_o;
reg hdmi2usbsoc_hdmi_in1_wer0_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_wer0_toggle_o;
reg hdmi2usbsoc_hdmi_in1_wer0_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_decoding0_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in1_decoding0_input;
reg hdmi2usbsoc_hdmi_in1_decoding0_valid_o = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_decoding0_output_raw = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_decoding0_output_d = 8'd0;
reg [1:0] hdmi2usbsoc_hdmi_in1_decoding0_output_c = 2'd0;
reg hdmi2usbsoc_hdmi_in1_decoding0_output_de = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_serdesstrobe;
reg [9:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_d = 10'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re;
wire [5:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r;
reg [5:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_w = 6'd0;
wire [1:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_busy_status;
wire [1:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_status;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_reset_re;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_reset_r;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_reset_w = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_se;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_delayed_master;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_delayed_slave;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_inc;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_ce;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_cal;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_rst;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_busy;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_cal;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_rst;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_busy;
wire [4:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr2;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_valid;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_incdec;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_edge;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_cascade;
reg [7:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness = 8'd128;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_too_late;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_too_early;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_reset_lateness;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_o_r = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_charsync1_raw_data;
reg hdmi2usbsoc_hdmi_in1_charsync1_synced = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_charsync1_data = 10'd0;
wire hdmi2usbsoc_hdmi_in1_charsync1_char_synced_status;
wire [3:0] hdmi2usbsoc_hdmi_in1_charsync1_ctl_pos_status;
reg [9:0] hdmi2usbsoc_hdmi_in1_charsync1_raw_data1 = 10'd0;
wire [19:0] hdmi2usbsoc_hdmi_in1_charsync1_raw;
reg hdmi2usbsoc_hdmi_in1_charsync1_found_control = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync1_control_position = 4'd0;
reg [2:0] hdmi2usbsoc_hdmi_in1_charsync1_control_counter = 3'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync1_previous_control_position = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync1_word_sel = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_wer1_data;
wire hdmi2usbsoc_hdmi_in1_wer1_update_re;
wire hdmi2usbsoc_hdmi_in1_wer1_update_r;
reg hdmi2usbsoc_hdmi_in1_wer1_update_w = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer1_status = 24'd0;
reg [8:0] hdmi2usbsoc_hdmi_in1_wer1_data_r = 9'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_wer1_transitions = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_wer1_transition_count = 4'd0;
reg hdmi2usbsoc_hdmi_in1_wer1_is_control = 1'd0;
reg hdmi2usbsoc_hdmi_in1_wer1_is_error = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer1_period_counter = 24'd0;
reg hdmi2usbsoc_hdmi_in1_wer1_period_done = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer1_wer_counter = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r = 24'd0;
reg hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r_updated = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer1_wer_counter_sys = 24'd0;
wire hdmi2usbsoc_hdmi_in1_wer1_i;
wire hdmi2usbsoc_hdmi_in1_wer1_o;
reg hdmi2usbsoc_hdmi_in1_wer1_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_wer1_toggle_o;
reg hdmi2usbsoc_hdmi_in1_wer1_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_decoding1_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in1_decoding1_input;
reg hdmi2usbsoc_hdmi_in1_decoding1_valid_o = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_decoding1_output_raw = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_decoding1_output_d = 8'd0;
reg [1:0] hdmi2usbsoc_hdmi_in1_decoding1_output_c = 2'd0;
reg hdmi2usbsoc_hdmi_in1_decoding1_output_de = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_serdesstrobe;
reg [9:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_d = 10'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re;
wire [5:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r;
reg [5:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_w = 6'd0;
wire [1:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_busy_status;
wire [1:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_status;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_reset_re;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_reset_r;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_reset_w = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_se;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_delayed_master;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_delayed_slave;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_inc;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_ce;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_cal;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_rst;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_busy;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_cal;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_rst;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_busy;
wire [4:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr2;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_valid;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_incdec;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_edge;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_cascade;
reg [7:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness = 8'd128;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_too_late;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_too_early;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_reset_lateness;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_master_pending = 1'd0;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_slave_pending = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_i;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_o;
reg hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_o_r = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_charsync2_raw_data;
reg hdmi2usbsoc_hdmi_in1_charsync2_synced = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_charsync2_data = 10'd0;
wire hdmi2usbsoc_hdmi_in1_charsync2_char_synced_status;
wire [3:0] hdmi2usbsoc_hdmi_in1_charsync2_ctl_pos_status;
reg [9:0] hdmi2usbsoc_hdmi_in1_charsync2_raw_data1 = 10'd0;
wire [19:0] hdmi2usbsoc_hdmi_in1_charsync2_raw;
reg hdmi2usbsoc_hdmi_in1_charsync2_found_control = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync2_control_position = 4'd0;
reg [2:0] hdmi2usbsoc_hdmi_in1_charsync2_control_counter = 3'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync2_previous_control_position = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_charsync2_word_sel = 4'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_wer2_data;
wire hdmi2usbsoc_hdmi_in1_wer2_update_re;
wire hdmi2usbsoc_hdmi_in1_wer2_update_r;
reg hdmi2usbsoc_hdmi_in1_wer2_update_w = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer2_status = 24'd0;
reg [8:0] hdmi2usbsoc_hdmi_in1_wer2_data_r = 9'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_wer2_transitions = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_wer2_transition_count = 4'd0;
reg hdmi2usbsoc_hdmi_in1_wer2_is_control = 1'd0;
reg hdmi2usbsoc_hdmi_in1_wer2_is_error = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer2_period_counter = 24'd0;
reg hdmi2usbsoc_hdmi_in1_wer2_period_done = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer2_wer_counter = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r = 24'd0;
reg hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r_updated = 1'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_wer2_wer_counter_sys = 24'd0;
wire hdmi2usbsoc_hdmi_in1_wer2_i;
wire hdmi2usbsoc_hdmi_in1_wer2_o;
reg hdmi2usbsoc_hdmi_in1_wer2_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_wer2_toggle_o;
reg hdmi2usbsoc_hdmi_in1_wer2_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_decoding2_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in1_decoding2_input;
reg hdmi2usbsoc_hdmi_in1_decoding2_valid_o = 1'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_decoding2_output_raw = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_decoding2_output_d = 8'd0;
reg [1:0] hdmi2usbsoc_hdmi_in1_decoding2_output_c = 2'd0;
reg hdmi2usbsoc_hdmi_in1_decoding2_output_de = 1'd0;
wire hdmi2usbsoc_hdmi_in1_chansync_valid_i;
reg hdmi2usbsoc_hdmi_in1_chansync_chan_synced = 1'd0;
wire hdmi2usbsoc_hdmi_in1_chansync_status;
wire hdmi2usbsoc_hdmi_in1_chansync_all_control;
wire [9:0] hdmi2usbsoc_hdmi_in1_chansync_data_in0_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_chansync_data_in0_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_chansync_data_in0_c;
wire hdmi2usbsoc_hdmi_in1_chansync_data_in0_de;
wire [9:0] hdmi2usbsoc_hdmi_in1_chansync_data_out0_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_chansync_data_out0_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_chansync_data_out0_c;
wire hdmi2usbsoc_hdmi_in1_chansync_data_out0_de;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_din;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_dout;
wire hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_re;
reg [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_produce = 3'd0;
reg [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_consume = 3'd0;
wire [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_we;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_w;
wire [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_rdport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in1_chansync_is_control0;
wire [9:0] hdmi2usbsoc_hdmi_in1_chansync_data_in1_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_chansync_data_in1_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_chansync_data_in1_c;
wire hdmi2usbsoc_hdmi_in1_chansync_data_in1_de;
wire [9:0] hdmi2usbsoc_hdmi_in1_chansync_data_out1_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_chansync_data_out1_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_chansync_data_out1_c;
wire hdmi2usbsoc_hdmi_in1_chansync_data_out1_de;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_din;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_dout;
wire hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_re;
reg [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_produce = 3'd0;
reg [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_consume = 3'd0;
wire [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_we;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_w;
wire [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_rdport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in1_chansync_is_control1;
wire [9:0] hdmi2usbsoc_hdmi_in1_chansync_data_in2_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_chansync_data_in2_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_chansync_data_in2_c;
wire hdmi2usbsoc_hdmi_in1_chansync_data_in2_de;
wire [9:0] hdmi2usbsoc_hdmi_in1_chansync_data_out2_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_chansync_data_out2_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_chansync_data_out2_c;
wire hdmi2usbsoc_hdmi_in1_chansync_data_out2_de;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_din;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_dout;
wire hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_re;
reg [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_produce = 3'd0;
reg [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_consume = 3'd0;
wire [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_we;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_w;
wire [2:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_rdport_adr;
wire [20:0] hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in1_chansync_is_control2;
wire hdmi2usbsoc_hdmi_in1_chansync_some_control;
wire hdmi2usbsoc_hdmi_in1_syncpol_valid_i;
wire [9:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in0_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in0_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in0_c;
wire hdmi2usbsoc_hdmi_in1_syncpol_data_in0_de;
wire [9:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in1_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in1_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in1_c;
wire hdmi2usbsoc_hdmi_in1_syncpol_data_in1_de;
wire [9:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in2_raw;
wire [7:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in2_d;
wire [1:0] hdmi2usbsoc_hdmi_in1_syncpol_data_in2_c;
wire hdmi2usbsoc_hdmi_in1_syncpol_data_in2_de;
reg hdmi2usbsoc_hdmi_in1_syncpol_valid_o = 1'd0;
wire hdmi2usbsoc_hdmi_in1_syncpol_de;
wire hdmi2usbsoc_hdmi_in1_syncpol_hsync;
wire hdmi2usbsoc_hdmi_in1_syncpol_vsync;
reg [7:0] hdmi2usbsoc_hdmi_in1_syncpol_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_syncpol_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_syncpol_b = 8'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_syncpol_c0 = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_syncpol_c1 = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_syncpol_c2 = 10'd0;
reg hdmi2usbsoc_hdmi_in1_syncpol_de_r = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_in1_syncpol_c_polarity = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_in1_syncpol_c_out = 2'd0;
wire hdmi2usbsoc_hdmi_in1_resdetection_valid_i;
wire hdmi2usbsoc_hdmi_in1_resdetection_vsync;
wire hdmi2usbsoc_hdmi_in1_resdetection_de;
wire [10:0] hdmi2usbsoc_hdmi_in1_resdetection_hres_status;
wire [10:0] hdmi2usbsoc_hdmi_in1_resdetection_vres_status;
reg hdmi2usbsoc_hdmi_in1_resdetection_de_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_resdetection_pn_de;
reg [10:0] hdmi2usbsoc_hdmi_in1_resdetection_hcounter = 11'd0;
reg [10:0] hdmi2usbsoc_hdmi_in1_resdetection_hcounter_st = 11'd0;
reg hdmi2usbsoc_hdmi_in1_resdetection_vsync_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_resdetection_p_vsync;
reg [10:0] hdmi2usbsoc_hdmi_in1_resdetection_vcounter = 11'd0;
reg [10:0] hdmi2usbsoc_hdmi_in1_resdetection_vcounter_st = 11'd0;
wire hdmi2usbsoc_hdmi_in1_frame_valid_i;
wire hdmi2usbsoc_hdmi_in1_frame_vsync;
wire hdmi2usbsoc_hdmi_in1_frame_de;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_r;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_g;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_b;
wire hdmi2usbsoc_hdmi_in1_frame_frame_valid;
wire hdmi2usbsoc_hdmi_in1_frame_frame_ready;
wire hdmi2usbsoc_hdmi_in1_frame_frame_first;
wire hdmi2usbsoc_hdmi_in1_frame_frame_last;
wire hdmi2usbsoc_hdmi_in1_frame_frame_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in1_frame_frame_payload_pixels;
wire hdmi2usbsoc_hdmi_in1_frame_busy;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_re;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_r;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_w;
reg hdmi2usbsoc_hdmi_in1_frame_de_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_valid;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_ready;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_last = 1'd0;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_b;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_valid;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_ready;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_first;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_last;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_cr;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_r;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_g;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_b;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_b = 8'd0;
reg signed [8:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_g = 9'sd0;
reg signed [8:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_g = 9'sd0;
reg signed [16:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_ca_mult_rg = 17'sd0;
reg signed [16:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb_mult_bg = 17'sd0;
reg signed [24:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_carg_plus_cbbg = 25'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw = 11'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_yraw = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_yraw = 12'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r0 = 11'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cc_mult_ryraw = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cd_mult_byraw = 20'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r1 = 11'sd0;
reg signed [10:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_y = 11'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cr = 12'sd0;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_ce;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce;
wire hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_busy;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n4 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n5 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n6 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n7 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n4 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n4 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n5 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n5 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n6 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n6 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n7 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n7 = 1'd0;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_valid;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_ready;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_first;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_cr;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_valid;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_ready;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_first;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_last;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_payload_cb_cr;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_y;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cb;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cr;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_cb_cr = 8'd0;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_cr = 8'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_parity = 1'd0;
reg [8:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cb_sum = 9'd0;
reg [8:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cr_sum = 9'd0;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cb_mean;
wire [7:0] hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cr_mean;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_ce;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce;
wire hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_busy;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync0 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync1 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync2 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de3 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync3 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de4 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync4 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de5 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync5 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de6 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync6 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de7 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync7 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de8 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync8 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de9 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync9 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_de10 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_next_vsync10 = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_vsync_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_frame_new_frame;
reg [63:0] hdmi2usbsoc_hdmi_in1_frame_cur_word = 64'd0;
reg hdmi2usbsoc_hdmi_in1_frame_cur_word_valid = 1'd0;
wire [15:0] hdmi2usbsoc_hdmi_in1_frame_encoded_pixel;
reg [1:0] hdmi2usbsoc_hdmi_in1_frame_pack_counter = 2'd0;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_sink_valid;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_in1_frame_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_fifo_sink_last = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_sof = 1'd0;
wire [63:0] hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_pixels;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_source_valid;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_source_ready;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_source_first;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_source_last;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_source_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in1_frame_fifo_source_payload_pixels;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_we;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_writable;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_re;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_readable;
wire [66:0] hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_din;
wire [66:0] hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_dout;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_ce;
(* register_balancing = "no" *) reg [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next;
reg [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_binary = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next_binary = 10'd0;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_ce;
(* register_balancing = "no" *) reg [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next;
reg [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_binary = 10'd0;
reg [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_produce_rdomain;
wire [9:0] hdmi2usbsoc_hdmi_in1_frame_fifo_consume_wdomain;
wire [8:0] hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_adr;
wire [66:0] hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_we;
wire [66:0] hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_dat_w;
wire [8:0] hdmi2usbsoc_hdmi_in1_frame_fifo_rdport_adr;
wire [66:0] hdmi2usbsoc_hdmi_in1_frame_fifo_rdport_dat_r;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_payload_pixels;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_last;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_payload_pixels;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_in1_frame_pix_overflow = 1'd0;
wire hdmi2usbsoc_hdmi_in1_frame_pix_overflow_reset;
wire hdmi2usbsoc_hdmi_in1_frame_sys_overflow;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_reset_i;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_reset_o;
reg hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_o;
reg hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_i;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_o;
reg hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_o;
reg hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_o_r = 1'd0;
reg hdmi2usbsoc_hdmi_in1_frame_overflow_mask = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_frame_valid;
reg hdmi2usbsoc_hdmi_in1_dma_frame_ready = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_frame_first;
wire hdmi2usbsoc_hdmi_in1_dma_frame_last;
wire hdmi2usbsoc_hdmi_in1_dma_frame_payload_sof;
wire [63:0] hdmi2usbsoc_hdmi_in1_dma_frame_payload_pixels;
reg [26:0] hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full = 27'd0;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_frame_size_storage;
reg hdmi2usbsoc_hdmi_in1_dma_frame_size_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_irq;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_address;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_address_reached;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_address_valid;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_address_done = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_pending;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_trigger;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_clear = 1'd0;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_reached;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_valid;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_done;
reg [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage_full = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_we;
wire [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_dat_w;
reg [26:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full = 27'd0;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_we;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_dat_w;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_pending;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_trigger;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_clear = 1'd0;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_reached;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_valid;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_done;
reg [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage_full = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_we;
wire [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_dat_w;
reg [26:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full = 27'd0;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_we;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_dat_w;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_status_re;
wire [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_status_r;
reg [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_status_w = 2'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_re;
wire [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_r;
reg [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_w = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_storage_full = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_in1_dma_slot_array_storage;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_re = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_slot_array_change_slot;
reg hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot = 1'd0;
reg hdmi2usbsoc_hdmi_in1_dma_reset_words = 1'd0;
reg hdmi2usbsoc_hdmi_in1_dma_count_word = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_last_word;
reg [23:0] hdmi2usbsoc_hdmi_in1_dma_current_address = 24'd0;
reg [23:0] hdmi2usbsoc_hdmi_in1_dma_mwords_remaining = 24'd0;
wire [63:0] hdmi2usbsoc_hdmi_in1_dma_memory_word;
reg hdmi2usbsoc_hdmi_in1_dma_sink_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_in1_dma_sink_sink_ready;
wire [23:0] hdmi2usbsoc_hdmi_in1_dma_sink_sink_payload_address;
wire [63:0] hdmi2usbsoc_hdmi_in1_dma_sink_sink_payload_data;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_sink_valid;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_in1_dma_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_in1_dma_fifo_sink_last = 1'd0;
wire [63:0] hdmi2usbsoc_hdmi_in1_dma_fifo_sink_payload_data;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_source_valid;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_source_ready;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_source_first;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_source_last;
wire [63:0] hdmi2usbsoc_hdmi_in1_dma_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_readable;
wire [65:0] hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_din;
wire [65:0] hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_dout;
reg [4:0] hdmi2usbsoc_hdmi_in1_dma_fifo_level = 5'd0;
reg hdmi2usbsoc_hdmi_in1_dma_fifo_replace = 1'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_dma_fifo_produce = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_dma_fifo_consume = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_adr = 4'd0;
wire [65:0] hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_we;
wire [65:0] hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_do_read;
wire [3:0] hdmi2usbsoc_hdmi_in1_dma_fifo_rdport_adr;
wire [65:0] hdmi2usbsoc_hdmi_in1_dma_fifo_rdport_dat_r;
wire [63:0] hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_last;
wire [63:0] hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_last;
wire hdmi2usbsoc_litedramport2_cmd_valid0;
wire hdmi2usbsoc_litedramport2_cmd_ready0;
wire hdmi2usbsoc_litedramport2_cmd_first0;
wire hdmi2usbsoc_litedramport2_cmd_last0;
wire hdmi2usbsoc_litedramport2_cmd_payload_we0;
wire [23:0] hdmi2usbsoc_litedramport2_cmd_payload_adr0;
wire hdmi2usbsoc_litedramport2_wdata_ready;
reg [63:0] hdmi2usbsoc_litedramport2_wdata_payload_data = 64'd0;
reg [7:0] hdmi2usbsoc_litedramport2_wdata_payload_we = 8'd0;
wire hdmi2usbsoc_litedramport2_rdata_valid0;
wire hdmi2usbsoc_litedramport2_rdata_ready0;
reg hdmi2usbsoc_litedramport2_rdata_first0 = 1'd0;
reg hdmi2usbsoc_litedramport2_rdata_last0 = 1'd0;
wire [63:0] hdmi2usbsoc_litedramport2_rdata_payload_data0;
reg hdmi2usbsoc_litedramport0_cmd_valid1 = 1'd0;
wire hdmi2usbsoc_litedramport0_cmd_ready1;
reg hdmi2usbsoc_litedramport0_cmd_first = 1'd0;
reg hdmi2usbsoc_litedramport0_cmd_last = 1'd0;
reg hdmi2usbsoc_litedramport0_cmd_payload_we1 = 1'd0;
reg [23:0] hdmi2usbsoc_litedramport0_cmd_payload_adr1 = 24'd0;
wire hdmi2usbsoc_litedramport0_rdata_valid1;
wire hdmi2usbsoc_litedramport0_rdata_ready;
wire hdmi2usbsoc_litedramport0_rdata_first;
wire hdmi2usbsoc_litedramport0_rdata_last;
wire [63:0] hdmi2usbsoc_litedramport0_rdata_payload_data1;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_valid;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_ready;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_first;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_last;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_payload_adr;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_valid;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_ready;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_first;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_last;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_payload_adr;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_we;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_writable;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_re;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_readable;
wire [26:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_din;
wire [26:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_dout;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_ce;
(* register_balancing = "no" *) reg [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q = 3'd0;
wire [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next;
reg [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_binary = 3'd0;
reg [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next_binary = 3'd0;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_ce;
(* register_balancing = "no" *) reg [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q = 3'd0;
wire [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next;
reg [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_binary = 3'd0;
reg [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary = 3'd0;
wire [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_produce_rdomain;
wire [2:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_consume_wdomain;
wire [1:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_adr;
wire [26:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_dat_r;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_we;
wire [26:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_dat_w;
wire [1:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_rdport_adr;
wire [26:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_rdport_dat_r;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_payload_adr;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_first;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_last;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_payload_adr;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_first;
wire hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_last;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_valid;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_ready;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_first;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_last;
wire [63:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_payload_data;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_valid;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_ready;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_first;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_last;
wire [63:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_payload_data;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_we;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_writable;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_re;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_readable;
wire [65:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_din;
wire [65:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_dout;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_ce;
(* register_balancing = "no" *) reg [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q = 5'd0;
wire [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next;
reg [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_binary = 5'd0;
reg [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next_binary = 5'd0;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_ce;
(* register_balancing = "no" *) reg [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q = 5'd0;
wire [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next;
reg [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_binary = 5'd0;
reg [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary = 5'd0;
wire [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_produce_rdomain;
wire [4:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_consume_wdomain;
wire [3:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_adr;
wire [65:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_dat_r;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_we;
wire [65:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_dat_w;
wire [3:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_rdport_adr;
wire [65:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_rdport_dat_r;
wire [63:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_first;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_last;
wire [63:0] hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_first;
wire hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_last;
wire hdmi2usbsoc_litedramport1_cmd_valid1;
reg hdmi2usbsoc_litedramport1_cmd_ready1 = 1'd0;
wire hdmi2usbsoc_litedramport1_cmd_payload_we1;
wire [25:0] hdmi2usbsoc_litedramport1_cmd_payload_adr1;
reg hdmi2usbsoc_litedramport1_rdata_valid1 = 1'd0;
wire hdmi2usbsoc_litedramport1_rdata_ready;
reg hdmi2usbsoc_litedramport1_rdata_first = 1'd0;
reg hdmi2usbsoc_litedramport1_rdata_last = 1'd0;
reg [15:0] hdmi2usbsoc_litedramport1_rdata_payload_data1 = 16'd0;
reg hdmi2usbsoc_litedramport1_flush = 1'd0;
reg hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_valid = 1'd0;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_ready;
reg hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_first = 1'd0;
reg hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_last = 1'd0;
reg [3:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_payload_sel = 4'd0;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_valid;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_ready;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_first;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_last;
wire [3:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_payload_sel;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_we;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_writable;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_re;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_readable;
wire [5:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_din;
wire [5:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_dout;
reg [2:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_level = 3'd0;
reg hdmi2usbsoc_litedramportconverter0_cmd_buffer_replace = 1'd0;
reg [1:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_produce = 2'd0;
reg [1:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_consume = 2'd0;
reg [1:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_adr = 2'd0;
wire [5:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_dat_r;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_we;
wire [5:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_dat_w;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_do_read;
wire [1:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_rdport_adr;
wire [5:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_rdport_dat_r;
wire [3:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_payload_sel;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_first;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_last;
wire [3:0] hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_payload_sel;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_first;
wire hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_last;
reg [1:0] hdmi2usbsoc_litedramportconverter0_counter = 2'd0;
reg hdmi2usbsoc_litedramportconverter0_counter_ce = 1'd0;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_valid;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_ready;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_last;
wire [63:0] hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_payload_data;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_valid;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_ready;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_last;
reg [63:0] hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_payload_data = 64'd0;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_pipe_ce;
wire hdmi2usbsoc_litedramportconverter0_rdata_buffer_busy;
reg hdmi2usbsoc_litedramportconverter0_rdata_buffer_valid_n = 1'd0;
reg hdmi2usbsoc_litedramportconverter0_rdata_buffer_first_n = 1'd0;
reg hdmi2usbsoc_litedramportconverter0_rdata_buffer_last_n = 1'd0;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_valid;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_ready;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_last;
wire [63:0] hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_payload_data;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_source_valid;
reg hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready = 1'd0;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_source_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_source_last;
wire [15:0] hdmi2usbsoc_litedramportconverter0_rdata_converter_source_payload_data;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_valid;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_ready;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_last;
reg [63:0] hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data = 64'd0;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_valid;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_ready;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_last;
reg [15:0] hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_data = 16'd0;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_valid_token_count;
reg [1:0] hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_mux = 2'd0;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_last;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_valid;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_ready;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_first;
wire hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_last;
wire [15:0] hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_payload_data;
reg [3:0] hdmi2usbsoc_litedramportconverter0_rdata_chunk = 4'd1;
wire hdmi2usbsoc_litedramportconverter0_rdata_chunk_valid;
wire hdmi2usbsoc_hdmi_out0_core_source_source_valid;
wire hdmi2usbsoc_hdmi_out0_core_source_source_ready;
wire [15:0] hdmi2usbsoc_hdmi_out0_core_source_source_payload_data;
wire hdmi2usbsoc_hdmi_out0_core_source_source_param_hsync;
wire hdmi2usbsoc_hdmi_out0_core_source_source_param_vsync;
wire hdmi2usbsoc_hdmi_out0_core_source_source_param_de;
reg hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage;
reg hdmi2usbsoc_hdmi_out0_core_underflow_enable_re = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_underflow_update_underflow_update_re;
wire hdmi2usbsoc_hdmi_out0_core_underflow_update_underflow_update_r;
reg hdmi2usbsoc_hdmi_out0_core_underflow_update_underflow_update_w = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi_out0_core_underflow_counter_status = 32'd0;
wire hdmi2usbsoc_hdmi_out0_core_initiator_source_source_valid;
wire hdmi2usbsoc_hdmi_out0_core_initiator_source_source_ready;
wire hdmi2usbsoc_hdmi_out0_core_initiator_source_source_first;
wire hdmi2usbsoc_hdmi_out0_core_initiator_source_source_last;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_length;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_valid;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_ready;
reg hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_last = 1'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_length;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_valid;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_ready;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_first;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_last;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_length;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_we;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_writable;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_re;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_readable;
wire [161:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_din;
wire [161:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_dout;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_ce;
(* register_balancing = "no" *) reg [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next;
reg [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary = 2'd0;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_ce;
(* register_balancing = "no" *) reg [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next;
reg [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_produce_rdomain;
wire [1:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_consume_wdomain;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_adr;
wire [161:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_we;
wire [161:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_rdport_adr;
wire [161:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_rdport_dat_r;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_length;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_first;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_last;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_length;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_first;
wire hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_last;
reg hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_enable_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_re = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_re = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage;
reg hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_re = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_valid;
wire hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_ready;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vscan;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_valid = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_ready = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_last = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_hsync = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_vsync = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_de = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_hactive = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_vactive = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_timinggenerator_active = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter = 12'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter = 12'd0;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_sink_valid;
reg hdmi2usbsoc_hdmi_out0_core_dmareader_sink_ready = 1'd0;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_dmareader_sink_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out0_core_dmareader_sink_payload_length;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_source_valid;
reg hdmi2usbsoc_hdmi_out0_core_dmareader_source_ready = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_source_first;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_source_last;
wire [15:0] hdmi2usbsoc_hdmi_out0_core_dmareader_source_payload_data;
reg hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_ready;
wire [25:0] hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_payload_address;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_valid;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_ready;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_first;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_last;
wire [15:0] hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_payload_data;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_request_enable;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_request_issued;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_data_dequeued;
reg [12:0] hdmi2usbsoc_hdmi_out0_core_dmareader_rsv_level = 13'd0;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_valid;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_ready;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_first;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_last;
wire [15:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_payload_data;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_first;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_last;
wire [15:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_re;
reg hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_readable = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_readable;
wire [17:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_din;
wire [17:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_dout;
reg [12:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 = 13'd0;
reg hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_replace = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_produce = 12'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_consume = 12'd0;
reg [11:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_adr = 12'd0;
wire [17:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_we;
wire [17:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_do_read;
wire [11:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_adr;
wire [17:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_dat_r;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_re;
wire [12:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level1;
wire [15:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_last;
wire [15:0] hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_last;
wire [25:0] hdmi2usbsoc_hdmi_out0_core_dmareader_base;
wire [25:0] hdmi2usbsoc_hdmi_out0_core_dmareader_length;
reg [25:0] hdmi2usbsoc_hdmi_out0_core_dmareader_offset = 26'd0;
wire hdmi2usbsoc_hdmi_out0_core_underflow_enable;
wire hdmi2usbsoc_hdmi_out0_core_underflow_update;
reg [31:0] hdmi2usbsoc_hdmi_out0_core_underflow_counter = 32'd0;
wire hdmi2usbsoc_hdmi_out0_core_i;
wire hdmi2usbsoc_hdmi_out0_core_o;
reg hdmi2usbsoc_hdmi_out0_core_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_out0_core_toggle_o;
reg hdmi2usbsoc_hdmi_out0_core_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_out0_driver_sink_sink_valid;
wire hdmi2usbsoc_hdmi_out0_driver_sink_sink_ready;
wire hdmi2usbsoc_hdmi_out0_driver_sink_sink_first;
wire hdmi2usbsoc_hdmi_out0_driver_sink_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_b;
wire hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_hsync;
wire hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_vsync;
wire hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_de;
reg [9:0] hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage_full = 10'd0;
wire [9:0] hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_re = 1'd0;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_re;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_r;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_w = 1'd0;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_send_go_re;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_send_go_r;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_send_go_w = 1'd0;
wire [3:0] hdmi2usbsoc_hdmi_out0_driver_clocking_status_status;
wire hdmi_out0_pix_clk;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_re = 1'd0;
reg [4:0] hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage_full = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_re = 1'd0;
wire [15:0] hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_r_status;
reg [15:0] hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage_full = 16'd0;
wire [15:0] hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_re = 1'd0;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_re;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_r;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_w = 1'd0;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_re;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_r;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_w = 1'd0;
reg hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy_status = 1'd0;
wire hdmi_out0_pix2x_clk;
wire hdmi_out0_pix10x_clk;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_serdesstrobe;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_clk_pix_unbuffered;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progdata;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progen;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progdone;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pix_locked;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_clocking_remaining_bits = 4'd0;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_transmitting;
reg [9:0] hdmi2usbsoc_hdmi_out0_driver_clocking_sr = 10'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_clocking_busy_counter = 4'd0;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_busy;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_mult_locked;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_clkfbout;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll_locked;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll0_pix10x;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll1_pix2x;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll2_pix;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_locked_async;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy;
wire hdmi2usbsoc_hdmi_out0_driver_clocking_hdmi_clk_se;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_valid;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_ready;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_first;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_b;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_hsync;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_vsync;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_de;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0;
wire [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_c;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_de;
reg [9:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1 = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1d = 4'd0;
reg [8:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m = 9'd0;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n;
reg [8:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r = 9'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m = 4'd0;
reg signed [5:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt = 6'sd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c0 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de0 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c1 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de1 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c2 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de2 = 1'd0;
reg [4:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x_pol = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_di;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_do;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_ti;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_to;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_pad_se;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0;
wire [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_c;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_de;
reg [9:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1 = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1d = 4'd0;
reg [8:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m = 9'd0;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n;
reg [8:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r = 9'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m = 4'd0;
reg signed [5:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt = 6'sd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c0 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de0 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c1 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de1 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c2 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de2 = 1'd0;
reg [4:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x_pol = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_di;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_do;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_ti;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_to;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_pad_se;
wire [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0;
wire [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_c;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_de;
reg [9:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1 = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1d = 4'd0;
reg [8:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m = 9'd0;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n;
reg [8:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r = 9'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m = 4'd0;
reg signed [5:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt = 6'sd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c0 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de0 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c1 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de1 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c2 = 2'd0;
reg hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de2 = 1'd0;
reg [4:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x_pol = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_di;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_do;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_ti;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_to;
wire hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_pad_se;
wire hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_valid;
reg hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready = 1'd0;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
wire hdmi2usbsoc_hdmi_out0_resetinserter_source_source_valid;
wire hdmi2usbsoc_hdmi_out0_resetinserter_source_source_ready;
reg hdmi2usbsoc_hdmi_out0_resetinserter_source_source_first = 1'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_source_source_last = 1'd0;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_cr;
reg hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_last = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_payload_data = 8'd0;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_dout;
reg [2:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level = 3'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_replace = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_produce = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_consume = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_do_read;
wire [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_last = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data = 8'd0;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_dout;
reg [2:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level = 3'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_replace = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_produce = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_consume = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_do_read;
wire [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_last = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data = 8'd0;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_dout;
reg [2:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level = 3'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_replace = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_produce = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_consume = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_do_read;
wire [1:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_out0_resetinserter_parity_in = 1'd0;
reg hdmi2usbsoc_hdmi_out0_resetinserter_parity_out = 1'd0;
wire hdmi2usbsoc_hdmi_out0_resetinserter_reset;
wire hdmi2usbsoc_hdmi_out0_sink_valid;
wire hdmi2usbsoc_hdmi_out0_sink_ready;
wire hdmi2usbsoc_hdmi_out0_sink_first;
wire hdmi2usbsoc_hdmi_out0_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_sink_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_out0_sink_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_out0_sink_payload_cr;
wire hdmi2usbsoc_hdmi_out0_source_valid;
wire hdmi2usbsoc_hdmi_out0_source_ready;
wire hdmi2usbsoc_hdmi_out0_source_first;
wire hdmi2usbsoc_hdmi_out0_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out0_source_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_out0_source_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_out0_source_payload_b;
wire [7:0] hdmi2usbsoc_hdmi_out0_sink_y;
wire [7:0] hdmi2usbsoc_hdmi_out0_sink_cb;
wire [7:0] hdmi2usbsoc_hdmi_out0_sink_cr;
reg [7:0] hdmi2usbsoc_hdmi_out0_source_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_source_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_source_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record3_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record3_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out0_record3_ycbcr_n_cr = 8'd0;
reg signed [8:0] hdmi2usbsoc_hdmi_out0_cb_minus_coffset = 9'sd0;
reg signed [8:0] hdmi2usbsoc_hdmi_out0_cr_minus_coffset = 9'sd0;
reg signed [8:0] hdmi2usbsoc_hdmi_out0_y_minus_yoffset = 9'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out0_cr_minus_coffset_mult_acoef = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out0_cb_minus_coffset_mult_bcoef = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out0_cr_minus_coffset_mult_ccoef = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out0_cb_minus_coffset_mult_dcoef = 20'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_out0_r = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_out0_g = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_out0_b = 12'sd0;
wire hdmi2usbsoc_hdmi_out0_ce;
wire hdmi2usbsoc_hdmi_out0_pipe_ce;
wire hdmi2usbsoc_hdmi_out0_busy;
reg hdmi2usbsoc_hdmi_out0_valid_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_valid_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_valid_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_valid_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_first_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_last_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_first_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_last_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_first_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_last_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_first_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_last_n3 = 1'd0;
wire hdmi2usbsoc_hdmi_out0_sink_payload_hsync;
wire hdmi2usbsoc_hdmi_out0_sink_payload_vsync;
wire hdmi2usbsoc_hdmi_out0_sink_payload_de;
wire hdmi2usbsoc_hdmi_out0_source_payload_hsync;
wire hdmi2usbsoc_hdmi_out0_source_payload_vsync;
wire hdmi2usbsoc_hdmi_out0_source_payload_de;
reg hdmi2usbsoc_hdmi_out0_next_s0 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s1 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s2 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s3 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s4 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s5 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s6 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s7 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s8 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s9 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s10 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s11 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s12 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s13 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s14 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s15 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s16 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_next_s17 = 1'd0;
reg hdmi2usbsoc_hdmi_out0_de_r = 1'd0;
reg hdmi2usbsoc_hdmi_out0_core_source_valid_d = 1'd0;
reg [15:0] hdmi2usbsoc_hdmi_out0_core_source_data_d = 16'd0;
wire hdmi2usbsoc_litedramport3_cmd_valid0;
wire hdmi2usbsoc_litedramport3_cmd_ready0;
wire hdmi2usbsoc_litedramport3_cmd_first;
wire hdmi2usbsoc_litedramport3_cmd_last;
wire hdmi2usbsoc_litedramport3_cmd_payload_we0;
wire [23:0] hdmi2usbsoc_litedramport3_cmd_payload_adr0;
wire hdmi2usbsoc_litedramport3_wdata_ready;
reg [63:0] hdmi2usbsoc_litedramport3_wdata_payload_data = 64'd0;
reg [7:0] hdmi2usbsoc_litedramport3_wdata_payload_we = 8'd0;
wire hdmi2usbsoc_litedramport3_rdata_valid0;
wire hdmi2usbsoc_litedramport3_rdata_ready0;
reg hdmi2usbsoc_litedramport3_rdata_first0 = 1'd0;
reg hdmi2usbsoc_litedramport3_rdata_last0 = 1'd0;
wire [63:0] hdmi2usbsoc_litedramport3_rdata_payload_data0;
reg hdmi2usbsoc_litedramport2_cmd_valid1 = 1'd0;
wire hdmi2usbsoc_litedramport2_cmd_ready1;
reg hdmi2usbsoc_litedramport2_cmd_first1 = 1'd0;
reg hdmi2usbsoc_litedramport2_cmd_last1 = 1'd0;
reg hdmi2usbsoc_litedramport2_cmd_payload_we1 = 1'd0;
reg [23:0] hdmi2usbsoc_litedramport2_cmd_payload_adr1 = 24'd0;
wire hdmi2usbsoc_litedramport2_rdata_valid1;
wire hdmi2usbsoc_litedramport2_rdata_ready1;
wire hdmi2usbsoc_litedramport2_rdata_first1;
wire hdmi2usbsoc_litedramport2_rdata_last1;
wire [63:0] hdmi2usbsoc_litedramport2_rdata_payload_data1;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_valid;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_ready;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_first;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_last;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_payload_adr;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_valid;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_ready;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_first;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_last;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_payload_adr;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_we;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_writable;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_re;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_readable;
wire [26:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_din;
wire [26:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_dout;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_ce;
(* register_balancing = "no" *) reg [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q = 3'd0;
wire [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next;
reg [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_binary = 3'd0;
reg [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next_binary = 3'd0;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_ce;
(* register_balancing = "no" *) reg [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q = 3'd0;
wire [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next;
reg [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_binary = 3'd0;
reg [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary = 3'd0;
wire [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_produce_rdomain;
wire [2:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_consume_wdomain;
wire [1:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_adr;
wire [26:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_dat_r;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_we;
wire [26:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_dat_w;
wire [1:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_rdport_adr;
wire [26:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_rdport_dat_r;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_payload_adr;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_first;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_last;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_payload_we;
wire [23:0] hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_payload_adr;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_first;
wire hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_last;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_valid;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_ready;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_first;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_last;
wire [63:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_payload_data;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_valid;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_ready;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_first;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_last;
wire [63:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_payload_data;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_we;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_writable;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_re;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_readable;
wire [65:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_din;
wire [65:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_dout;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_ce;
(* register_balancing = "no" *) reg [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q = 5'd0;
wire [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next;
reg [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_binary = 5'd0;
reg [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next_binary = 5'd0;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_ce;
(* register_balancing = "no" *) reg [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q = 5'd0;
wire [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next;
reg [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_binary = 5'd0;
reg [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary = 5'd0;
wire [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_produce_rdomain;
wire [4:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_consume_wdomain;
wire [3:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_adr;
wire [65:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_dat_r;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_we;
wire [65:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_dat_w;
wire [3:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_rdport_adr;
wire [65:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_rdport_dat_r;
wire [63:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_first;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_last;
wire [63:0] hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_first;
wire hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_last;
wire hdmi2usbsoc_litedramport3_cmd_valid1;
reg hdmi2usbsoc_litedramport3_cmd_ready1 = 1'd0;
wire hdmi2usbsoc_litedramport3_cmd_payload_we1;
wire [25:0] hdmi2usbsoc_litedramport3_cmd_payload_adr1;
reg hdmi2usbsoc_litedramport3_rdata_valid1 = 1'd0;
wire hdmi2usbsoc_litedramport3_rdata_ready1;
reg hdmi2usbsoc_litedramport3_rdata_first1 = 1'd0;
reg hdmi2usbsoc_litedramport3_rdata_last1 = 1'd0;
reg [15:0] hdmi2usbsoc_litedramport3_rdata_payload_data1 = 16'd0;
reg hdmi2usbsoc_litedramport3_flush = 1'd0;
reg hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_valid = 1'd0;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_ready;
reg hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_first = 1'd0;
reg hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_last = 1'd0;
reg [3:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_payload_sel = 4'd0;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_valid;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_ready;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_first;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_last;
wire [3:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_payload_sel;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_we;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_writable;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_re;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_readable;
wire [5:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_din;
wire [5:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_dout;
reg [2:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_level = 3'd0;
reg hdmi2usbsoc_litedramportconverter1_cmd_buffer_replace = 1'd0;
reg [1:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_produce = 2'd0;
reg [1:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_consume = 2'd0;
reg [1:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_adr = 2'd0;
wire [5:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_dat_r;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_we;
wire [5:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_dat_w;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_do_read;
wire [1:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_rdport_adr;
wire [5:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_rdport_dat_r;
wire [3:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_payload_sel;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_first;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_last;
wire [3:0] hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_payload_sel;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_first;
wire hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_last;
reg [1:0] hdmi2usbsoc_litedramportconverter1_counter = 2'd0;
reg hdmi2usbsoc_litedramportconverter1_counter_ce = 1'd0;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_valid;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_ready;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_last;
wire [63:0] hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_payload_data;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_valid;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_ready;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_last;
reg [63:0] hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_payload_data = 64'd0;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_pipe_ce;
wire hdmi2usbsoc_litedramportconverter1_rdata_buffer_busy;
reg hdmi2usbsoc_litedramportconverter1_rdata_buffer_valid_n = 1'd0;
reg hdmi2usbsoc_litedramportconverter1_rdata_buffer_first_n = 1'd0;
reg hdmi2usbsoc_litedramportconverter1_rdata_buffer_last_n = 1'd0;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_valid;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_ready;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_last;
wire [63:0] hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_payload_data;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_source_valid;
reg hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready = 1'd0;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_source_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_source_last;
wire [15:0] hdmi2usbsoc_litedramportconverter1_rdata_converter_source_payload_data;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_valid;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_ready;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_last;
reg [63:0] hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data = 64'd0;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_valid;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_ready;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_last;
reg [15:0] hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_data = 16'd0;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_valid_token_count;
reg [1:0] hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_mux = 2'd0;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_last;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_valid;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_ready;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_first;
wire hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_last;
wire [15:0] hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_payload_data;
reg [3:0] hdmi2usbsoc_litedramportconverter1_rdata_chunk = 4'd1;
wire hdmi2usbsoc_litedramportconverter1_rdata_chunk_valid;
wire hdmi2usbsoc_hdmi_out1_core_source_source_valid;
wire hdmi2usbsoc_hdmi_out1_core_source_source_ready;
wire [15:0] hdmi2usbsoc_hdmi_out1_core_source_source_payload_data;
wire hdmi2usbsoc_hdmi_out1_core_source_source_param_hsync;
wire hdmi2usbsoc_hdmi_out1_core_source_source_param_vsync;
wire hdmi2usbsoc_hdmi_out1_core_source_source_param_de;
reg hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage;
reg hdmi2usbsoc_hdmi_out1_core_underflow_enable_re = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_underflow_update_underflow_update_re;
wire hdmi2usbsoc_hdmi_out1_core_underflow_update_underflow_update_r;
reg hdmi2usbsoc_hdmi_out1_core_underflow_update_underflow_update_w = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi_out1_core_underflow_counter_status = 32'd0;
wire hdmi2usbsoc_hdmi_out1_core_initiator_source_source_valid;
wire hdmi2usbsoc_hdmi_out1_core_initiator_source_source_ready;
wire hdmi2usbsoc_hdmi_out1_core_initiator_source_source_first;
wire hdmi2usbsoc_hdmi_out1_core_initiator_source_source_last;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_length;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_valid;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_ready;
reg hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_last = 1'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_length;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_valid;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_ready;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_first;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_last;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_length;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_we;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_writable;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_re;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_readable;
wire [161:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_din;
wire [161:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_dout;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_ce;
(* register_balancing = "no" *) reg [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next;
reg [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_binary = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next_binary = 2'd0;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_ce;
(* register_balancing = "no" *) reg [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next;
reg [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_binary = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary = 2'd0;
wire [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_produce_rdomain;
wire [1:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_consume_wdomain;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_adr;
wire [161:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_we;
wire [161:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_rdport_adr;
wire [161:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_rdport_dat_r;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_length;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_first;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_last;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vscan;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_length;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_first;
wire hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_last;
reg hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage_full = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_enable_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_re = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage_full = 12'd0;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_re = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_re = 1'd0;
reg [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full = 32'd0;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage;
reg hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_re = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_valid;
wire hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_ready;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hscan;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vres;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vsync_start;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vsync_end;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vscan;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_valid = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_ready = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_last = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_hsync = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_vsync = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_de = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_hactive = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_vactive = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_timinggenerator_active = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter = 12'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter = 12'd0;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_sink_valid;
reg hdmi2usbsoc_hdmi_out1_core_dmareader_sink_ready = 1'd0;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_dmareader_sink_payload_base;
wire [31:0] hdmi2usbsoc_hdmi_out1_core_dmareader_sink_payload_length;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_source_valid;
reg hdmi2usbsoc_hdmi_out1_core_dmareader_source_ready = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_source_first;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_source_last;
wire [15:0] hdmi2usbsoc_hdmi_out1_core_dmareader_source_payload_data;
reg hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_ready;
wire [25:0] hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_payload_address;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_valid;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_ready;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_first;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_last;
wire [15:0] hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_payload_data;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_request_enable;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_request_issued;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_data_dequeued;
reg [12:0] hdmi2usbsoc_hdmi_out1_core_dmareader_rsv_level = 13'd0;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_valid;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_ready;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_first;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_last;
wire [15:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_payload_data;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_first;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_last;
wire [15:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_re;
reg hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_readable = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_readable;
wire [17:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_din;
wire [17:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_dout;
reg [12:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 = 13'd0;
reg hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_replace = 1'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_produce = 12'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_consume = 12'd0;
reg [11:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_adr = 12'd0;
wire [17:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_we;
wire [17:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_do_read;
wire [11:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_adr;
wire [17:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_dat_r;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_re;
wire [12:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level1;
wire [15:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_last;
wire [15:0] hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_last;
wire [25:0] hdmi2usbsoc_hdmi_out1_core_dmareader_base;
wire [25:0] hdmi2usbsoc_hdmi_out1_core_dmareader_length;
reg [25:0] hdmi2usbsoc_hdmi_out1_core_dmareader_offset = 26'd0;
wire hdmi2usbsoc_hdmi_out1_core_underflow_enable;
wire hdmi2usbsoc_hdmi_out1_core_underflow_update;
reg [31:0] hdmi2usbsoc_hdmi_out1_core_underflow_counter = 32'd0;
wire hdmi2usbsoc_hdmi_out1_core_i;
wire hdmi2usbsoc_hdmi_out1_core_o;
reg hdmi2usbsoc_hdmi_out1_core_toggle_i = 1'd0;
wire hdmi2usbsoc_hdmi_out1_core_toggle_o;
reg hdmi2usbsoc_hdmi_out1_core_toggle_o_r = 1'd0;
wire hdmi2usbsoc_hdmi_out1_driver_sink_sink_valid;
wire hdmi2usbsoc_hdmi_out1_driver_sink_sink_ready;
wire hdmi2usbsoc_hdmi_out1_driver_sink_sink_first;
wire hdmi2usbsoc_hdmi_out1_driver_sink_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_b;
wire hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_hsync;
wire hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_vsync;
wire hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_de;
wire hdmi_out1_pix_clk;
wire hdmi_out1_pix2x_clk;
wire hdmi_out1_pix10x_clk;
wire hdmi2usbsoc_hdmi_out1_driver_clocking_serdesstrobe;
wire hdmi2usbsoc_hdmi_out1_driver_clocking_hdmi_clk_se;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_valid;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_ready;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_first;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_b;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_hsync;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_vsync;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_de;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0;
wire [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_c;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_de;
reg [9:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1 = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1d = 4'd0;
reg [8:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m = 9'd0;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n;
reg [8:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r = 9'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m = 4'd0;
reg signed [5:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt = 6'sd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c0 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de0 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c1 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de1 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c2 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de2 = 1'd0;
reg [4:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x_pol = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_di;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_do;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_ti;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_to;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_pad_se;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0;
wire [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_c;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_de;
reg [9:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1 = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1d = 4'd0;
reg [8:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m = 9'd0;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n;
reg [8:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r = 9'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m = 4'd0;
reg signed [5:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt = 6'sd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c0 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de0 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c1 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de1 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c2 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de2 = 1'd0;
reg [4:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x_pol = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_di;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_do;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_ti;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_to;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_pad_se;
wire [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0;
wire [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_c;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_de;
reg [9:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out = 10'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1 = 8'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1d = 4'd0;
reg [8:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m = 9'd0;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n;
reg [8:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r = 9'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m = 4'd0;
reg [3:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m = 4'd0;
reg signed [5:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt = 6'sd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c0 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de0 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c1 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de1 = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c2 = 2'd0;
reg hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de2 = 1'd0;
reg [4:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x_pol = 5'd0;
wire [4:0] hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_di;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_do;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_ti;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_to;
wire hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_pad_se;
wire hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_valid;
reg hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready = 1'd0;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_cb_cr;
wire hdmi2usbsoc_hdmi_out1_resetinserter_source_source_valid;
wire hdmi2usbsoc_hdmi_out1_resetinserter_source_source_ready;
reg hdmi2usbsoc_hdmi_out1_resetinserter_source_source_first = 1'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_source_source_last = 1'd0;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_cr;
reg hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_last = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_payload_data = 8'd0;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_dout;
reg [2:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level = 3'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_replace = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_produce = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_consume = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_do_read;
wire [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_last = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_payload_data = 8'd0;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_dout;
reg [2:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level = 3'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_replace = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_produce = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_consume = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_do_read;
wire [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_valid = 1'd0;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_ready;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_first = 1'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_last = 1'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_payload_data = 8'd0;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_valid;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_ready;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_we;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_writable;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_re;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_readable;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_din;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_dout;
reg [2:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level = 3'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_replace = 1'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_produce = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_consume = 2'd0;
reg [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_adr = 2'd0;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_dat_r;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_we;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_dat_w;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_do_read;
wire [1:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_rdport_adr;
wire [9:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_rdport_dat_r;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_payload_data;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_first;
wire hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_last;
reg hdmi2usbsoc_hdmi_out1_resetinserter_parity_in = 1'd0;
reg hdmi2usbsoc_hdmi_out1_resetinserter_parity_out = 1'd0;
wire hdmi2usbsoc_hdmi_out1_resetinserter_reset;
wire hdmi2usbsoc_hdmi_out1_sink_valid;
wire hdmi2usbsoc_hdmi_out1_sink_ready;
wire hdmi2usbsoc_hdmi_out1_sink_first;
wire hdmi2usbsoc_hdmi_out1_sink_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_sink_payload_y;
wire [7:0] hdmi2usbsoc_hdmi_out1_sink_payload_cb;
wire [7:0] hdmi2usbsoc_hdmi_out1_sink_payload_cr;
wire hdmi2usbsoc_hdmi_out1_source_valid;
wire hdmi2usbsoc_hdmi_out1_source_ready;
wire hdmi2usbsoc_hdmi_out1_source_first;
wire hdmi2usbsoc_hdmi_out1_source_last;
wire [7:0] hdmi2usbsoc_hdmi_out1_source_payload_r;
wire [7:0] hdmi2usbsoc_hdmi_out1_source_payload_g;
wire [7:0] hdmi2usbsoc_hdmi_out1_source_payload_b;
wire [7:0] hdmi2usbsoc_hdmi_out1_sink_y;
wire [7:0] hdmi2usbsoc_hdmi_out1_sink_cb;
wire [7:0] hdmi2usbsoc_hdmi_out1_sink_cr;
reg [7:0] hdmi2usbsoc_hdmi_out1_source_r = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_source_g = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_source_b = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_cr = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record3_ycbcr_n_y = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record3_ycbcr_n_cb = 8'd0;
reg [7:0] hdmi2usbsoc_hdmi_out1_record3_ycbcr_n_cr = 8'd0;
reg signed [8:0] hdmi2usbsoc_hdmi_out1_cb_minus_coffset = 9'sd0;
reg signed [8:0] hdmi2usbsoc_hdmi_out1_cr_minus_coffset = 9'sd0;
reg signed [8:0] hdmi2usbsoc_hdmi_out1_y_minus_yoffset = 9'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out1_cr_minus_coffset_mult_acoef = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out1_cb_minus_coffset_mult_bcoef = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out1_cr_minus_coffset_mult_ccoef = 20'sd0;
reg signed [19:0] hdmi2usbsoc_hdmi_out1_cb_minus_coffset_mult_dcoef = 20'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_out1_r = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_out1_g = 12'sd0;
reg signed [11:0] hdmi2usbsoc_hdmi_out1_b = 12'sd0;
wire hdmi2usbsoc_hdmi_out1_ce;
wire hdmi2usbsoc_hdmi_out1_pipe_ce;
wire hdmi2usbsoc_hdmi_out1_busy;
reg hdmi2usbsoc_hdmi_out1_valid_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_valid_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_valid_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_valid_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_first_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_last_n0 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_first_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_last_n1 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_first_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_last_n2 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_first_n3 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_last_n3 = 1'd0;
wire hdmi2usbsoc_hdmi_out1_sink_payload_hsync;
wire hdmi2usbsoc_hdmi_out1_sink_payload_vsync;
wire hdmi2usbsoc_hdmi_out1_sink_payload_de;
wire hdmi2usbsoc_hdmi_out1_source_payload_hsync;
wire hdmi2usbsoc_hdmi_out1_source_payload_vsync;
wire hdmi2usbsoc_hdmi_out1_source_payload_de;
reg hdmi2usbsoc_hdmi_out1_next_s0 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s1 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s2 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s3 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s4 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s5 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s6 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s7 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s8 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s9 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s10 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s11 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s12 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s13 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s14 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s15 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s16 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_next_s17 = 1'd0;
reg hdmi2usbsoc_hdmi_out1_de_r = 1'd0;
reg hdmi2usbsoc_hdmi_out1_core_source_valid_d = 1'd0;
reg [15:0] hdmi2usbsoc_hdmi_out1_core_source_data_d = 16'd0;
reg encoder_port_port_cmd_valid = 1'd0;
wire encoder_port_port_cmd_ready;
reg encoder_port_port_cmd_payload_we = 1'd0;
reg [23:0] encoder_port_port_cmd_payload_adr = 24'd0;
wire encoder_port_port_wdata_ready;
reg [63:0] encoder_port_port_wdata_payload_data = 64'd0;
reg [7:0] encoder_port_port_wdata_payload_we = 8'd0;
wire encoder_port_port_rdata_valid;
wire encoder_port_port_rdata_ready;
reg encoder_port_port_rdata_first = 1'd0;
reg encoder_port_port_rdata_last = 1'd0;
wire [63:0] encoder_port_port_rdata_payload_data;
wire encoder_port_new_port_cmd_valid;
reg encoder_port_new_port_cmd_ready = 1'd0;
wire encoder_port_new_port_cmd_payload_we;
wire [22:0] encoder_port_new_port_cmd_payload_adr;
wire encoder_port_new_port_rdata_valid;
wire encoder_port_new_port_rdata_ready;
wire encoder_port_new_port_rdata_first;
wire encoder_port_new_port_rdata_last;
wire [127:0] encoder_port_new_port_rdata_payload_data;
reg encoder_port_counter = 1'd0;
reg encoder_port_counter_reset = 1'd0;
reg encoder_port_counter_ce = 1'd0;
wire encoder_port_sink_valid;
wire encoder_port_sink_ready;
wire encoder_port_sink_first;
wire encoder_port_sink_last;
wire [63:0] encoder_port_sink_payload_data;
wire encoder_port_source_valid;
wire encoder_port_source_ready;
wire encoder_port_source_first;
wire encoder_port_source_last;
reg [127:0] encoder_port_source_payload_data = 128'd0;
wire encoder_port_converter_sink_valid;
wire encoder_port_converter_sink_ready;
wire encoder_port_converter_sink_first;
wire encoder_port_converter_sink_last;
wire [63:0] encoder_port_converter_sink_payload_data;
wire encoder_port_converter_source_valid;
wire encoder_port_converter_source_ready;
reg encoder_port_converter_source_first = 1'd0;
reg encoder_port_converter_source_last = 1'd0;
reg [127:0] encoder_port_converter_source_payload_data = 128'd0;
reg [1:0] encoder_port_converter_source_payload_valid_token_count = 2'd0;
reg encoder_port_converter_demux = 1'd0;
wire encoder_port_converter_load_part;
reg encoder_port_converter_strobe_all = 1'd0;
wire encoder_port_source_source_valid;
wire encoder_port_source_source_ready;
wire encoder_port_source_source_first;
wire encoder_port_source_source_last;
wire [127:0] encoder_port_source_source_payload_data;
wire encoder_reader_source_valid;
wire encoder_reader_source_ready;
wire encoder_reader_source_first;
wire encoder_reader_source_last;
wire [127:0] encoder_reader_source_payload_data;
reg [31:0] encoder_reader_base_storage_full = 32'd0;
wire [31:0] encoder_reader_base_storage;
reg encoder_reader_base_re = 1'd0;
reg [15:0] encoder_reader_h_width_storage_full = 16'd0;
wire [15:0] encoder_reader_h_width_storage;
reg encoder_reader_h_width_re = 1'd0;
reg [15:0] encoder_reader_v_width_storage_full = 16'd0;
wire [15:0] encoder_reader_v_width_storage;
reg encoder_reader_v_width_re = 1'd0;
wire encoder_reader_start_re;
wire encoder_reader_start_r;
reg encoder_reader_start_w = 1'd0;
reg encoder_reader_status = 1'd0;
reg encoder_reader_sink_sink_valid = 1'd0;
wire encoder_reader_sink_sink_ready;
wire [22:0] encoder_reader_sink_sink_payload_address;
wire encoder_reader_source_source_valid;
wire encoder_reader_source_source_ready;
wire encoder_reader_source_source_first;
wire encoder_reader_source_source_last;
wire [127:0] encoder_reader_source_source_payload_data;
wire encoder_reader_request_enable;
wire encoder_reader_request_issued;
wire encoder_reader_data_dequeued;
reg [4:0] encoder_reader_rsv_level = 5'd0;
wire encoder_reader_fifo_sink_valid;
wire encoder_reader_fifo_sink_ready;
wire encoder_reader_fifo_sink_first;
wire encoder_reader_fifo_sink_last;
wire [127:0] encoder_reader_fifo_sink_payload_data;
wire encoder_reader_fifo_source_valid;
wire encoder_reader_fifo_source_ready;
wire encoder_reader_fifo_source_first;
wire encoder_reader_fifo_source_last;
wire [127:0] encoder_reader_fifo_source_payload_data;
wire encoder_reader_fifo_syncfifo_we;
wire encoder_reader_fifo_syncfifo_writable;
wire encoder_reader_fifo_syncfifo_re;
wire encoder_reader_fifo_syncfifo_readable;
wire [129:0] encoder_reader_fifo_syncfifo_din;
wire [129:0] encoder_reader_fifo_syncfifo_dout;
reg [4:0] encoder_reader_fifo_level = 5'd0;
reg encoder_reader_fifo_replace = 1'd0;
reg [3:0] encoder_reader_fifo_produce = 4'd0;
reg [3:0] encoder_reader_fifo_consume = 4'd0;
reg [3:0] encoder_reader_fifo_wrport_adr = 4'd0;
wire [129:0] encoder_reader_fifo_wrport_dat_r;
wire encoder_reader_fifo_wrport_we;
wire [129:0] encoder_reader_fifo_wrport_dat_w;
wire encoder_reader_fifo_do_read;
wire [3:0] encoder_reader_fifo_rdport_adr;
wire [129:0] encoder_reader_fifo_rdport_dat_r;
wire [127:0] encoder_reader_fifo_fifo_in_payload_data;
wire encoder_reader_fifo_fifo_in_first;
wire encoder_reader_fifo_fifo_in_last;
wire [127:0] encoder_reader_fifo_fifo_out_payload_data;
wire encoder_reader_fifo_fifo_out_first;
wire encoder_reader_fifo_fifo_out_last;
reg [31:0] encoder_reader_base = 32'd0;
reg encoder_reader_h_clr = 1'd0;
reg encoder_reader_h_clr_lsb = 1'd0;
reg encoder_reader_h_inc = 1'd0;
reg [15:0] encoder_reader_h = 16'd0;
wire [15:0] encoder_reader_h_next;
reg encoder_reader_v_clr = 1'd0;
reg encoder_reader_v_inc = 1'd0;
reg encoder_reader_v_dec7 = 1'd0;
reg [15:0] encoder_reader_v = 16'd0;
wire [26:0] encoder_reader_read_address;
wire encoder_cdc_sink_valid;
wire encoder_cdc_sink_ready;
wire encoder_cdc_sink_first;
wire encoder_cdc_sink_last;
wire [127:0] encoder_cdc_sink_payload_data;
wire encoder_cdc_source_valid;
wire encoder_cdc_source_ready;
wire encoder_cdc_source_first;
wire encoder_cdc_source_last;
wire [127:0] encoder_cdc_source_payload_data;
wire encoder_cdc_asyncfifo_we;
wire encoder_cdc_asyncfifo_writable;
wire encoder_cdc_asyncfifo_re;
wire encoder_cdc_asyncfifo_readable;
wire [129:0] encoder_cdc_asyncfifo_din;
wire [129:0] encoder_cdc_asyncfifo_dout;
wire encoder_cdc_graycounter0_ce;
(* register_balancing = "no" *) reg [2:0] encoder_cdc_graycounter0_q = 3'd0;
wire [2:0] encoder_cdc_graycounter0_q_next;
reg [2:0] encoder_cdc_graycounter0_q_binary = 3'd0;
reg [2:0] encoder_cdc_graycounter0_q_next_binary = 3'd0;
wire encoder_cdc_graycounter1_ce;
(* register_balancing = "no" *) reg [2:0] encoder_cdc_graycounter1_q = 3'd0;
wire [2:0] encoder_cdc_graycounter1_q_next;
reg [2:0] encoder_cdc_graycounter1_q_binary = 3'd0;
reg [2:0] encoder_cdc_graycounter1_q_next_binary = 3'd0;
wire [2:0] encoder_cdc_produce_rdomain;
wire [2:0] encoder_cdc_consume_wdomain;
wire [1:0] encoder_cdc_wrport_adr;
wire [129:0] encoder_cdc_wrport_dat_r;
wire encoder_cdc_wrport_we;
wire [129:0] encoder_cdc_wrport_dat_w;
wire [1:0] encoder_cdc_rdport_adr;
wire [129:0] encoder_cdc_rdport_dat_r;
wire [127:0] encoder_cdc_fifo_in_payload_data;
wire encoder_cdc_fifo_in_first;
wire encoder_cdc_fifo_in_last;
wire [127:0] encoder_cdc_fifo_out_payload_data;
wire encoder_cdc_fifo_out_first;
wire encoder_cdc_fifo_out_last;
wire encoderbuffer_sink_valid;
reg encoderbuffer_sink_ready = 1'd0;
wire encoderbuffer_sink_first;
wire encoderbuffer_sink_last;
wire [127:0] encoderbuffer_sink_payload_data;
reg encoderbuffer_source_valid = 1'd0;
wire encoderbuffer_source_ready;
reg encoderbuffer_source_first = 1'd0;
reg encoderbuffer_source_last = 1'd0;
reg [15:0] encoderbuffer_source_payload_data = 16'd0;
reg [3:0] encoderbuffer_write_port_adr = 4'd0;
wire [127:0] encoderbuffer_write_port_dat_r;
wire encoderbuffer_write_port_we;
wire [127:0] encoderbuffer_write_port_dat_w;
reg [3:0] encoderbuffer_read_port_adr = 4'd0;
wire [127:0] encoderbuffer_read_port_dat_r;
reg encoderbuffer_write_sel = 1'd0;
reg encoderbuffer_write_swap = 1'd0;
reg encoderbuffer_read_sel = 1'd1;
reg encoderbuffer_read_swap = 1'd0;
reg encoderbuffer_v_write_clr = 1'd0;
reg encoderbuffer_v_write_inc = 1'd0;
reg [2:0] encoderbuffer_v_write = 3'd0;
reg encoderbuffer_h_read_clr = 1'd0;
reg encoderbuffer_h_read_inc = 1'd0;
reg [2:0] encoderbuffer_h_read = 3'd0;
reg encoderbuffer_v_read_clr = 1'd0;
reg encoderbuffer_v_read_inc = 1'd0;
reg [2:0] encoderbuffer_v_read = 3'd0;
wire encoder_sink_sink_valid0;
wire encoder_sink_sink_ready0;
wire encoder_sink_sink_first0;
wire encoder_sink_sink_last0;
wire [15:0] encoder_sink_sink_payload_data;
wire encoder_source_source_valid0;
wire encoder_source_source_ready0;
wire encoder_source_source_first;
wire encoder_source_source_last;
wire [7:0] encoder_source_source_payload_data;
wire [29:0] encoder_bus_adr;
wire [31:0] encoder_bus_dat_w;
wire [31:0] encoder_bus_dat_r;
wire [3:0] encoder_bus_sel;
wire encoder_bus_cyc;
wire encoder_bus_stb;
wire encoder_bus_ack;
wire encoder_bus_we;
wire [2:0] encoder_bus_cti;
wire [1:0] encoder_bus_bte;
wire encoder_bus_err;
wire encoder_sink_sink_valid1;
reg encoder_sink_sink_ready1 = 1'd0;
wire encoder_sink_sink_first1;
wire encoder_sink_sink_last1;
wire [7:0] encoder_sink_sink_payload_y;
wire [7:0] encoder_sink_sink_payload_cb_cr;
wire encoder_source_source_valid1;
wire encoder_source_source_ready1;
wire [7:0] encoder_source_source_payload_y;
wire [7:0] encoder_source_source_payload_cb;
wire [7:0] encoder_source_source_payload_cr;
reg encoder_y_fifo_sink_valid = 1'd0;
wire encoder_y_fifo_sink_ready;
reg encoder_y_fifo_sink_first = 1'd0;
reg encoder_y_fifo_sink_last = 1'd0;
reg [7:0] encoder_y_fifo_sink_payload_data = 8'd0;
wire encoder_y_fifo_source_valid;
wire encoder_y_fifo_source_ready;
wire encoder_y_fifo_source_first;
wire encoder_y_fifo_source_last;
wire [7:0] encoder_y_fifo_source_payload_data;
wire encoder_y_fifo_syncfifo_we;
wire encoder_y_fifo_syncfifo_writable;
wire encoder_y_fifo_syncfifo_re;
wire encoder_y_fifo_syncfifo_readable;
wire [9:0] encoder_y_fifo_syncfifo_din;
wire [9:0] encoder_y_fifo_syncfifo_dout;
reg [2:0] encoder_y_fifo_level = 3'd0;
reg encoder_y_fifo_replace = 1'd0;
reg [1:0] encoder_y_fifo_produce = 2'd0;
reg [1:0] encoder_y_fifo_consume = 2'd0;
reg [1:0] encoder_y_fifo_wrport_adr = 2'd0;
wire [9:0] encoder_y_fifo_wrport_dat_r;
wire encoder_y_fifo_wrport_we;
wire [9:0] encoder_y_fifo_wrport_dat_w;
wire encoder_y_fifo_do_read;
wire [1:0] encoder_y_fifo_rdport_adr;
wire [9:0] encoder_y_fifo_rdport_dat_r;
wire [7:0] encoder_y_fifo_fifo_in_payload_data;
wire encoder_y_fifo_fifo_in_first;
wire encoder_y_fifo_fifo_in_last;
wire [7:0] encoder_y_fifo_fifo_out_payload_data;
wire encoder_y_fifo_fifo_out_first;
wire encoder_y_fifo_fifo_out_last;
reg encoder_cb_fifo_sink_valid = 1'd0;
wire encoder_cb_fifo_sink_ready;
reg encoder_cb_fifo_sink_first = 1'd0;
reg encoder_cb_fifo_sink_last = 1'd0;
reg [7:0] encoder_cb_fifo_sink_payload_data = 8'd0;
wire encoder_cb_fifo_source_valid;
wire encoder_cb_fifo_source_ready;
wire encoder_cb_fifo_source_first;
wire encoder_cb_fifo_source_last;
wire [7:0] encoder_cb_fifo_source_payload_data;
wire encoder_cb_fifo_syncfifo_we;
wire encoder_cb_fifo_syncfifo_writable;
wire encoder_cb_fifo_syncfifo_re;
wire encoder_cb_fifo_syncfifo_readable;
wire [9:0] encoder_cb_fifo_syncfifo_din;
wire [9:0] encoder_cb_fifo_syncfifo_dout;
reg [2:0] encoder_cb_fifo_level = 3'd0;
reg encoder_cb_fifo_replace = 1'd0;
reg [1:0] encoder_cb_fifo_produce = 2'd0;
reg [1:0] encoder_cb_fifo_consume = 2'd0;
reg [1:0] encoder_cb_fifo_wrport_adr = 2'd0;
wire [9:0] encoder_cb_fifo_wrport_dat_r;
wire encoder_cb_fifo_wrport_we;
wire [9:0] encoder_cb_fifo_wrport_dat_w;
wire encoder_cb_fifo_do_read;
wire [1:0] encoder_cb_fifo_rdport_adr;
wire [9:0] encoder_cb_fifo_rdport_dat_r;
wire [7:0] encoder_cb_fifo_fifo_in_payload_data;
wire encoder_cb_fifo_fifo_in_first;
wire encoder_cb_fifo_fifo_in_last;
wire [7:0] encoder_cb_fifo_fifo_out_payload_data;
wire encoder_cb_fifo_fifo_out_first;
wire encoder_cb_fifo_fifo_out_last;
reg encoder_cr_fifo_sink_valid = 1'd0;
wire encoder_cr_fifo_sink_ready;
reg encoder_cr_fifo_sink_first = 1'd0;
reg encoder_cr_fifo_sink_last = 1'd0;
reg [7:0] encoder_cr_fifo_sink_payload_data = 8'd0;
wire encoder_cr_fifo_source_valid;
wire encoder_cr_fifo_source_ready;
wire encoder_cr_fifo_source_first;
wire encoder_cr_fifo_source_last;
wire [7:0] encoder_cr_fifo_source_payload_data;
wire encoder_cr_fifo_syncfifo_we;
wire encoder_cr_fifo_syncfifo_writable;
wire encoder_cr_fifo_syncfifo_re;
wire encoder_cr_fifo_syncfifo_readable;
wire [9:0] encoder_cr_fifo_syncfifo_din;
wire [9:0] encoder_cr_fifo_syncfifo_dout;
reg [2:0] encoder_cr_fifo_level = 3'd0;
reg encoder_cr_fifo_replace = 1'd0;
reg [1:0] encoder_cr_fifo_produce = 2'd0;
reg [1:0] encoder_cr_fifo_consume = 2'd0;
reg [1:0] encoder_cr_fifo_wrport_adr = 2'd0;
wire [9:0] encoder_cr_fifo_wrport_dat_r;
wire encoder_cr_fifo_wrport_we;
wire [9:0] encoder_cr_fifo_wrport_dat_w;
wire encoder_cr_fifo_do_read;
wire [1:0] encoder_cr_fifo_rdport_adr;
wire [9:0] encoder_cr_fifo_rdport_dat_r;
wire [7:0] encoder_cr_fifo_fifo_in_payload_data;
wire encoder_cr_fifo_fifo_in_first;
wire encoder_cr_fifo_fifo_in_last;
wire [7:0] encoder_cr_fifo_fifo_out_payload_data;
wire encoder_cr_fifo_fifo_out_first;
wire encoder_cr_fifo_fifo_out_last;
reg encoder_parity_in = 1'd0;
reg encoder_parity_out = 1'd0;
reg encoder_reset = 1'd0;
wire encoder_fdct_fifo_rd;
wire [23:0] encoder_fdct_fifo_q;
wire encoder_fdct_fifo_hf_full;
reg [23:0] encoder_fdct_data_d1 = 24'd0;
reg [23:0] encoder_fdct_data_d2 = 24'd0;
reg [23:0] encoder_fdct_data_d3 = 24'd0;
reg [23:0] encoder_fdct_data_d4 = 24'd0;
reg [23:0] encoder_fdct_data_d5 = 24'd0;
wire encoder_output_fifo_almost_full;
wire encoder_output_fifo_sink_valid;
wire encoder_output_fifo_sink_ready;
reg encoder_output_fifo_sink_first = 1'd0;
reg encoder_output_fifo_sink_last = 1'd0;
wire [7:0] encoder_output_fifo_sink_payload_data;
wire encoder_output_fifo_source_valid;
wire encoder_output_fifo_source_ready;
wire encoder_output_fifo_source_first;
wire encoder_output_fifo_source_last;
wire [7:0] encoder_output_fifo_source_payload_data;
wire encoder_output_fifo_re;
reg encoder_output_fifo_readable = 1'd0;
wire encoder_output_fifo_syncfifo_we;
wire encoder_output_fifo_syncfifo_writable;
wire encoder_output_fifo_syncfifo_re;
wire encoder_output_fifo_syncfifo_readable;
wire [9:0] encoder_output_fifo_syncfifo_din;
wire [9:0] encoder_output_fifo_syncfifo_dout;
reg [10:0] encoder_output_fifo_level0 = 11'd0;
reg encoder_output_fifo_replace = 1'd0;
reg [9:0] encoder_output_fifo_produce = 10'd0;
reg [9:0] encoder_output_fifo_consume = 10'd0;
reg [9:0] encoder_output_fifo_wrport_adr = 10'd0;
wire [9:0] encoder_output_fifo_wrport_dat_r;
wire encoder_output_fifo_wrport_we;
wire [9:0] encoder_output_fifo_wrport_dat_w;
wire encoder_output_fifo_do_read;
wire [9:0] encoder_output_fifo_rdport_adr;
wire [9:0] encoder_output_fifo_rdport_dat_r;
wire encoder_output_fifo_rdport_re;
wire [10:0] encoder_output_fifo_level1;
wire [7:0] encoder_output_fifo_fifo_in_payload_data;
wire encoder_output_fifo_fifo_in_first;
wire encoder_output_fifo_fifo_in_last;
wire [7:0] encoder_output_fifo_fifo_out_payload_data;
wire encoder_output_fifo_fifo_out_first;
wire encoder_output_fifo_fifo_out_last;
wire [29:0] encoder_jpeg_bus_adr;
wire [31:0] encoder_jpeg_bus_dat_w;
wire [31:0] encoder_jpeg_bus_dat_r;
wire [3:0] encoder_jpeg_bus_sel;
wire encoder_jpeg_bus_cyc;
wire encoder_jpeg_bus_stb;
wire encoder_jpeg_bus_ack;
wire encoder_jpeg_bus_we;
wire encoder_jpeg_bus_err;
reg [1:0] encoder = 2'd0;
wire encoder_streamer_sink_sink_valid;
wire encoder_streamer_sink_sink_ready;
wire encoder_streamer_sink_sink_first;
wire encoder_streamer_sink_sink_last;
wire [7:0] encoder_streamer_sink_sink_payload_data;
(* keep = "true" *) wire usb_clk;
wire usb_rst;
wire encoder_streamer_fifo_sink_valid;
wire encoder_streamer_fifo_sink_ready;
wire encoder_streamer_fifo_sink_first;
wire encoder_streamer_fifo_sink_last;
wire [7:0] encoder_streamer_fifo_sink_payload_data;
wire encoder_streamer_fifo_source_valid;
wire encoder_streamer_fifo_source_ready;
wire encoder_streamer_fifo_source_first;
wire encoder_streamer_fifo_source_last;
wire [7:0] encoder_streamer_fifo_source_payload_data;
wire encoder_streamer_fifo_asyncfifo_we;
wire encoder_streamer_fifo_asyncfifo_writable;
wire encoder_streamer_fifo_asyncfifo_re;
wire encoder_streamer_fifo_asyncfifo_readable;
wire [9:0] encoder_streamer_fifo_asyncfifo_din;
wire [9:0] encoder_streamer_fifo_asyncfifo_dout;
wire encoder_streamer_fifo_graycounter0_ce;
(* register_balancing = "no" *) reg [2:0] encoder_streamer_fifo_graycounter0_q = 3'd0;
wire [2:0] encoder_streamer_fifo_graycounter0_q_next;
reg [2:0] encoder_streamer_fifo_graycounter0_q_binary = 3'd0;
reg [2:0] encoder_streamer_fifo_graycounter0_q_next_binary = 3'd0;
wire encoder_streamer_fifo_graycounter1_ce;
(* register_balancing = "no" *) reg [2:0] encoder_streamer_fifo_graycounter1_q = 3'd0;
wire [2:0] encoder_streamer_fifo_graycounter1_q_next;
reg [2:0] encoder_streamer_fifo_graycounter1_q_binary = 3'd0;
reg [2:0] encoder_streamer_fifo_graycounter1_q_next_binary = 3'd0;
wire [2:0] encoder_streamer_fifo_produce_rdomain;
wire [2:0] encoder_streamer_fifo_consume_wdomain;
wire [1:0] encoder_streamer_fifo_wrport_adr;
wire [9:0] encoder_streamer_fifo_wrport_dat_r;
wire encoder_streamer_fifo_wrport_we;
wire [9:0] encoder_streamer_fifo_wrport_dat_w;
wire [1:0] encoder_streamer_fifo_rdport_adr;
wire [9:0] encoder_streamer_fifo_rdport_dat_r;
wire [7:0] encoder_streamer_fifo_fifo_in_payload_data;
wire encoder_streamer_fifo_fifo_in_first;
wire encoder_streamer_fifo_fifo_in_last;
wire [7:0] encoder_streamer_fifo_fifo_out_payload_data;
wire encoder_streamer_fifo_fifo_out_first;
wire encoder_streamer_fifo_fifo_out_last;
reg [1:0] controllerinjector_refresher_state = 2'd0;
reg [1:0] controllerinjector_refresher_next_state = 2'd0;
reg [2:0] controllerinjector_bankmachine0_state = 3'd0;
reg [2:0] controllerinjector_bankmachine0_next_state = 3'd0;
reg [2:0] controllerinjector_bankmachine1_state = 3'd0;
reg [2:0] controllerinjector_bankmachine1_next_state = 3'd0;
reg [2:0] controllerinjector_bankmachine2_state = 3'd0;
reg [2:0] controllerinjector_bankmachine2_next_state = 3'd0;
reg [2:0] controllerinjector_bankmachine3_state = 3'd0;
reg [2:0] controllerinjector_bankmachine3_next_state = 3'd0;
reg [2:0] controllerinjector_bankmachine4_state = 3'd0;
reg [2:0] controllerinjector_bankmachine4_next_state = 3'd0;
reg [2:0] controllerinjector_bankmachine5_state = 3'd0;
reg [2:0] controllerinjector_bankmachine5_next_state = 3'd0;
reg [2:0] controllerinjector_bankmachine6_state = 3'd0;
reg [2:0] controllerinjector_bankmachine6_next_state = 3'd0;
reg [2:0] controllerinjector_bankmachine7_state = 3'd0;
reg [2:0] controllerinjector_bankmachine7_next_state = 3'd0;
reg [3:0] controllerinjector_multiplexer_state = 4'd0;
reg [3:0] controllerinjector_multiplexer_next_state = 4'd0;
reg controllerinjector_state = 1'd0;
reg controllerinjector_next_state = 1'd0;
wire [2:0] controllerinjector_cba0;
wire [20:0] controllerinjector_rca0;
wire [2:0] controllerinjector_cba1;
wire [20:0] controllerinjector_rca1;
wire [2:0] controllerinjector_cba2;
wire [20:0] controllerinjector_rca2;
wire [2:0] controllerinjector_cba3;
wire [20:0] controllerinjector_rca3;
wire [2:0] controllerinjector_cba4;
wire [20:0] controllerinjector_rca4;
wire [2:0] controllerinjector_cba5;
wire [20:0] controllerinjector_rca5;
wire [5:0] controllerinjector_roundrobin0_request;
reg [2:0] controllerinjector_roundrobin0_grant = 3'd0;
wire controllerinjector_roundrobin0_ce;
wire [5:0] controllerinjector_roundrobin1_request;
reg [2:0] controllerinjector_roundrobin1_grant = 3'd0;
wire controllerinjector_roundrobin1_ce;
wire [5:0] controllerinjector_roundrobin2_request;
reg [2:0] controllerinjector_roundrobin2_grant = 3'd0;
wire controllerinjector_roundrobin2_ce;
wire [5:0] controllerinjector_roundrobin3_request;
reg [2:0] controllerinjector_roundrobin3_grant = 3'd0;
wire controllerinjector_roundrobin3_ce;
wire [5:0] controllerinjector_roundrobin4_request;
reg [2:0] controllerinjector_roundrobin4_grant = 3'd0;
wire controllerinjector_roundrobin4_ce;
wire [5:0] controllerinjector_roundrobin5_request;
reg [2:0] controllerinjector_roundrobin5_grant = 3'd0;
wire controllerinjector_roundrobin5_ce;
wire [5:0] controllerinjector_roundrobin6_request;
reg [2:0] controllerinjector_roundrobin6_grant = 3'd0;
wire controllerinjector_roundrobin6_ce;
wire [5:0] controllerinjector_roundrobin7_request;
reg [2:0] controllerinjector_roundrobin7_grant = 3'd0;
wire controllerinjector_roundrobin7_ce;
reg controllerinjector_new_master_wdata_ready0 = 1'd0;
reg controllerinjector_new_master_wdata_ready1 = 1'd0;
reg controllerinjector_new_master_wdata_ready2 = 1'd0;
reg controllerinjector_new_master_wdata_ready3 = 1'd0;
reg controllerinjector_new_master_wdata_ready4 = 1'd0;
reg controllerinjector_new_master_wdata_ready5 = 1'd0;
reg controllerinjector_new_master_rdata_valid0 = 1'd0;
reg controllerinjector_new_master_rdata_valid1 = 1'd0;
reg controllerinjector_new_master_rdata_valid2 = 1'd0;
reg controllerinjector_new_master_rdata_valid3 = 1'd0;
reg controllerinjector_new_master_rdata_valid4 = 1'd0;
reg controllerinjector_new_master_rdata_valid5 = 1'd0;
reg controllerinjector_new_master_rdata_valid6 = 1'd0;
reg controllerinjector_new_master_rdata_valid7 = 1'd0;
reg controllerinjector_new_master_rdata_valid8 = 1'd0;
reg controllerinjector_new_master_rdata_valid9 = 1'd0;
reg controllerinjector_new_master_rdata_valid10 = 1'd0;
reg controllerinjector_new_master_rdata_valid11 = 1'd0;
reg controllerinjector_new_master_rdata_valid12 = 1'd0;
reg controllerinjector_new_master_rdata_valid13 = 1'd0;
reg controllerinjector_new_master_rdata_valid14 = 1'd0;
reg controllerinjector_new_master_rdata_valid15 = 1'd0;
reg controllerinjector_new_master_rdata_valid16 = 1'd0;
reg controllerinjector_new_master_rdata_valid17 = 1'd0;
reg controllerinjector_new_master_rdata_valid18 = 1'd0;
reg controllerinjector_new_master_rdata_valid19 = 1'd0;
reg controllerinjector_new_master_rdata_valid20 = 1'd0;
reg controllerinjector_new_master_rdata_valid21 = 1'd0;
reg controllerinjector_new_master_rdata_valid22 = 1'd0;
reg controllerinjector_new_master_rdata_valid23 = 1'd0;
reg controllerinjector_new_master_rdata_valid24 = 1'd0;
reg controllerinjector_new_master_rdata_valid25 = 1'd0;
reg controllerinjector_new_master_rdata_valid26 = 1'd0;
reg controllerinjector_new_master_rdata_valid27 = 1'd0;
reg controllerinjector_new_master_rdata_valid28 = 1'd0;
reg controllerinjector_new_master_rdata_valid29 = 1'd0;
reg controllerinjector_new_master_rdata_valid30 = 1'd0;
reg controllerinjector_new_master_rdata_valid31 = 1'd0;
reg controllerinjector_new_master_rdata_valid32 = 1'd0;
reg controllerinjector_new_master_rdata_valid33 = 1'd0;
reg controllerinjector_new_master_rdata_valid34 = 1'd0;
reg controllerinjector_new_master_rdata_valid35 = 1'd0;
reg [2:0] cache_state = 3'd0;
reg [2:0] cache_next_state = 3'd0;
reg [1:0] litedramwishbonebridge_state = 2'd0;
reg [1:0] litedramwishbonebridge_next_state = 2'd0;
reg [3:0] edid0_state = 4'd0;
reg [3:0] edid0_next_state = 4'd0;
reg [1:0] dma0_state = 2'd0;
reg [1:0] dma0_next_state = 2'd0;
reg [3:0] edid1_state = 4'd0;
reg [3:0] edid1_next_state = 4'd0;
reg [1:0] dma1_state = 2'd0;
reg [1:0] dma1_next_state = 2'd0;
reg videoout0_state = 1'd0;
reg videoout0_next_state = 1'd0;
reg [25:0] hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value = 26'd0;
reg hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value_ce = 1'd0;
reg videoout1_state = 1'd0;
reg videoout1_next_state = 1'd0;
reg [25:0] hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value = 26'd0;
reg hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value_ce = 1'd0;
reg encoderdmareader_state = 1'd0;
reg encoderdmareader_next_state = 1'd0;
reg fsm0_state = 1'd0;
reg fsm0_next_state = 1'd0;
reg fsm1_state = 1'd0;
reg fsm1_next_state = 1'd0;
wire wb_sdram_con_request;
wire wb_sdram_con_grant;
wire [29:0] hdmi2usbsoc_shared_adr;
wire [31:0] hdmi2usbsoc_shared_dat_w;
wire [31:0] hdmi2usbsoc_shared_dat_r;
wire [3:0] hdmi2usbsoc_shared_sel;
wire hdmi2usbsoc_shared_cyc;
wire hdmi2usbsoc_shared_stb;
wire hdmi2usbsoc_shared_ack;
wire hdmi2usbsoc_shared_we;
wire [2:0] hdmi2usbsoc_shared_cti;
wire [1:0] hdmi2usbsoc_shared_bte;
wire hdmi2usbsoc_shared_err;
wire [1:0] hdmi2usbsoc_request;
reg hdmi2usbsoc_grant = 1'd0;
reg [5:0] hdmi2usbsoc_slave_sel = 6'd0;
reg [5:0] hdmi2usbsoc_slave_sel_r = 6'd0;
wire [13:0] hdmi2usbsoc_interface0_bank_bus_adr;
wire hdmi2usbsoc_interface0_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface0_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface0_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank0_base3_re;
wire [7:0] hdmi2usbsoc_csrbank0_base3_r;
wire [7:0] hdmi2usbsoc_csrbank0_base3_w;
wire hdmi2usbsoc_csrbank0_base2_re;
wire [7:0] hdmi2usbsoc_csrbank0_base2_r;
wire [7:0] hdmi2usbsoc_csrbank0_base2_w;
wire hdmi2usbsoc_csrbank0_base1_re;
wire [7:0] hdmi2usbsoc_csrbank0_base1_r;
wire [7:0] hdmi2usbsoc_csrbank0_base1_w;
wire hdmi2usbsoc_csrbank0_base0_re;
wire [7:0] hdmi2usbsoc_csrbank0_base0_r;
wire [7:0] hdmi2usbsoc_csrbank0_base0_w;
wire hdmi2usbsoc_csrbank0_h_width1_re;
wire [7:0] hdmi2usbsoc_csrbank0_h_width1_r;
wire [7:0] hdmi2usbsoc_csrbank0_h_width1_w;
wire hdmi2usbsoc_csrbank0_h_width0_re;
wire [7:0] hdmi2usbsoc_csrbank0_h_width0_r;
wire [7:0] hdmi2usbsoc_csrbank0_h_width0_w;
wire hdmi2usbsoc_csrbank0_v_width1_re;
wire [7:0] hdmi2usbsoc_csrbank0_v_width1_r;
wire [7:0] hdmi2usbsoc_csrbank0_v_width1_w;
wire hdmi2usbsoc_csrbank0_v_width0_re;
wire [7:0] hdmi2usbsoc_csrbank0_v_width0_r;
wire [7:0] hdmi2usbsoc_csrbank0_v_width0_w;
wire hdmi2usbsoc_csrbank0_done_re;
wire hdmi2usbsoc_csrbank0_done_r;
wire hdmi2usbsoc_csrbank0_done_w;
wire hdmi2usbsoc_csrbank0_sel;
wire [13:0] hdmi2usbsoc_interface0_sram_bus_adr;
wire hdmi2usbsoc_interface0_sram_bus_we;
wire [7:0] hdmi2usbsoc_interface0_sram_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface0_sram_bus_dat_r = 8'd0;
wire [6:0] hdmi2usbsoc_sram0_adr;
wire [7:0] hdmi2usbsoc_sram0_dat_r;
wire hdmi2usbsoc_sram0_we;
wire [7:0] hdmi2usbsoc_sram0_dat_w;
wire hdmi2usbsoc_sram0_sel;
reg hdmi2usbsoc_sram0_sel_r = 1'd0;
wire [13:0] hdmi2usbsoc_interface1_bank_bus_adr;
wire hdmi2usbsoc_interface1_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface1_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface1_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank1_edid_hpd_notif_re;
wire hdmi2usbsoc_csrbank1_edid_hpd_notif_r;
wire hdmi2usbsoc_csrbank1_edid_hpd_notif_w;
wire hdmi2usbsoc_csrbank1_edid_hpd_en0_re;
wire hdmi2usbsoc_csrbank1_edid_hpd_en0_r;
wire hdmi2usbsoc_csrbank1_edid_hpd_en0_w;
wire hdmi2usbsoc_csrbank1_clocking_pll_reset0_re;
wire hdmi2usbsoc_csrbank1_clocking_pll_reset0_r;
wire hdmi2usbsoc_csrbank1_clocking_pll_reset0_w;
wire hdmi2usbsoc_csrbank1_clocking_locked_re;
wire hdmi2usbsoc_csrbank1_clocking_locked_r;
wire hdmi2usbsoc_csrbank1_clocking_locked_w;
wire hdmi2usbsoc_csrbank1_clocking_pll_adr0_re;
wire [4:0] hdmi2usbsoc_csrbank1_clocking_pll_adr0_r;
wire [4:0] hdmi2usbsoc_csrbank1_clocking_pll_adr0_w;
wire hdmi2usbsoc_csrbank1_clocking_pll_dat_r1_re;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_r1_r;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_r1_w;
wire hdmi2usbsoc_csrbank1_clocking_pll_dat_r0_re;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_r0_r;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_r0_w;
wire hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_re;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_r;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_w;
wire hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_re;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_r;
wire [7:0] hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_w;
wire hdmi2usbsoc_csrbank1_clocking_pll_drdy_re;
wire hdmi2usbsoc_csrbank1_clocking_pll_drdy_r;
wire hdmi2usbsoc_csrbank1_clocking_pll_drdy_w;
wire hdmi2usbsoc_csrbank1_data0_cap_dly_busy_re;
wire [1:0] hdmi2usbsoc_csrbank1_data0_cap_dly_busy_r;
wire [1:0] hdmi2usbsoc_csrbank1_data0_cap_dly_busy_w;
wire hdmi2usbsoc_csrbank1_data0_cap_phase_re;
wire [1:0] hdmi2usbsoc_csrbank1_data0_cap_phase_r;
wire [1:0] hdmi2usbsoc_csrbank1_data0_cap_phase_w;
wire hdmi2usbsoc_csrbank1_data0_charsync_char_synced_re;
wire hdmi2usbsoc_csrbank1_data0_charsync_char_synced_r;
wire hdmi2usbsoc_csrbank1_data0_charsync_char_synced_w;
wire hdmi2usbsoc_csrbank1_data0_charsync_ctl_pos_re;
wire [3:0] hdmi2usbsoc_csrbank1_data0_charsync_ctl_pos_r;
wire [3:0] hdmi2usbsoc_csrbank1_data0_charsync_ctl_pos_w;
wire hdmi2usbsoc_csrbank1_data0_wer_value2_re;
wire [7:0] hdmi2usbsoc_csrbank1_data0_wer_value2_r;
wire [7:0] hdmi2usbsoc_csrbank1_data0_wer_value2_w;
wire hdmi2usbsoc_csrbank1_data0_wer_value1_re;
wire [7:0] hdmi2usbsoc_csrbank1_data0_wer_value1_r;
wire [7:0] hdmi2usbsoc_csrbank1_data0_wer_value1_w;
wire hdmi2usbsoc_csrbank1_data0_wer_value0_re;
wire [7:0] hdmi2usbsoc_csrbank1_data0_wer_value0_r;
wire [7:0] hdmi2usbsoc_csrbank1_data0_wer_value0_w;
wire hdmi2usbsoc_csrbank1_data1_cap_dly_busy_re;
wire [1:0] hdmi2usbsoc_csrbank1_data1_cap_dly_busy_r;
wire [1:0] hdmi2usbsoc_csrbank1_data1_cap_dly_busy_w;
wire hdmi2usbsoc_csrbank1_data1_cap_phase_re;
wire [1:0] hdmi2usbsoc_csrbank1_data1_cap_phase_r;
wire [1:0] hdmi2usbsoc_csrbank1_data1_cap_phase_w;
wire hdmi2usbsoc_csrbank1_data1_charsync_char_synced_re;
wire hdmi2usbsoc_csrbank1_data1_charsync_char_synced_r;
wire hdmi2usbsoc_csrbank1_data1_charsync_char_synced_w;
wire hdmi2usbsoc_csrbank1_data1_charsync_ctl_pos_re;
wire [3:0] hdmi2usbsoc_csrbank1_data1_charsync_ctl_pos_r;
wire [3:0] hdmi2usbsoc_csrbank1_data1_charsync_ctl_pos_w;
wire hdmi2usbsoc_csrbank1_data1_wer_value2_re;
wire [7:0] hdmi2usbsoc_csrbank1_data1_wer_value2_r;
wire [7:0] hdmi2usbsoc_csrbank1_data1_wer_value2_w;
wire hdmi2usbsoc_csrbank1_data1_wer_value1_re;
wire [7:0] hdmi2usbsoc_csrbank1_data1_wer_value1_r;
wire [7:0] hdmi2usbsoc_csrbank1_data1_wer_value1_w;
wire hdmi2usbsoc_csrbank1_data1_wer_value0_re;
wire [7:0] hdmi2usbsoc_csrbank1_data1_wer_value0_r;
wire [7:0] hdmi2usbsoc_csrbank1_data1_wer_value0_w;
wire hdmi2usbsoc_csrbank1_data2_cap_dly_busy_re;
wire [1:0] hdmi2usbsoc_csrbank1_data2_cap_dly_busy_r;
wire [1:0] hdmi2usbsoc_csrbank1_data2_cap_dly_busy_w;
wire hdmi2usbsoc_csrbank1_data2_cap_phase_re;
wire [1:0] hdmi2usbsoc_csrbank1_data2_cap_phase_r;
wire [1:0] hdmi2usbsoc_csrbank1_data2_cap_phase_w;
wire hdmi2usbsoc_csrbank1_data2_charsync_char_synced_re;
wire hdmi2usbsoc_csrbank1_data2_charsync_char_synced_r;
wire hdmi2usbsoc_csrbank1_data2_charsync_char_synced_w;
wire hdmi2usbsoc_csrbank1_data2_charsync_ctl_pos_re;
wire [3:0] hdmi2usbsoc_csrbank1_data2_charsync_ctl_pos_r;
wire [3:0] hdmi2usbsoc_csrbank1_data2_charsync_ctl_pos_w;
wire hdmi2usbsoc_csrbank1_data2_wer_value2_re;
wire [7:0] hdmi2usbsoc_csrbank1_data2_wer_value2_r;
wire [7:0] hdmi2usbsoc_csrbank1_data2_wer_value2_w;
wire hdmi2usbsoc_csrbank1_data2_wer_value1_re;
wire [7:0] hdmi2usbsoc_csrbank1_data2_wer_value1_r;
wire [7:0] hdmi2usbsoc_csrbank1_data2_wer_value1_w;
wire hdmi2usbsoc_csrbank1_data2_wer_value0_re;
wire [7:0] hdmi2usbsoc_csrbank1_data2_wer_value0_r;
wire [7:0] hdmi2usbsoc_csrbank1_data2_wer_value0_w;
wire hdmi2usbsoc_csrbank1_chansync_channels_synced_re;
wire hdmi2usbsoc_csrbank1_chansync_channels_synced_r;
wire hdmi2usbsoc_csrbank1_chansync_channels_synced_w;
wire hdmi2usbsoc_csrbank1_resdetection_hres1_re;
wire [2:0] hdmi2usbsoc_csrbank1_resdetection_hres1_r;
wire [2:0] hdmi2usbsoc_csrbank1_resdetection_hres1_w;
wire hdmi2usbsoc_csrbank1_resdetection_hres0_re;
wire [7:0] hdmi2usbsoc_csrbank1_resdetection_hres0_r;
wire [7:0] hdmi2usbsoc_csrbank1_resdetection_hres0_w;
wire hdmi2usbsoc_csrbank1_resdetection_vres1_re;
wire [2:0] hdmi2usbsoc_csrbank1_resdetection_vres1_r;
wire [2:0] hdmi2usbsoc_csrbank1_resdetection_vres1_w;
wire hdmi2usbsoc_csrbank1_resdetection_vres0_re;
wire [7:0] hdmi2usbsoc_csrbank1_resdetection_vres0_r;
wire [7:0] hdmi2usbsoc_csrbank1_resdetection_vres0_w;
wire hdmi2usbsoc_csrbank1_dma_frame_size3_re;
wire [2:0] hdmi2usbsoc_csrbank1_dma_frame_size3_r;
wire [2:0] hdmi2usbsoc_csrbank1_dma_frame_size3_w;
wire hdmi2usbsoc_csrbank1_dma_frame_size2_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_frame_size2_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_frame_size2_w;
wire hdmi2usbsoc_csrbank1_dma_frame_size1_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_frame_size1_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_frame_size1_w;
wire hdmi2usbsoc_csrbank1_dma_frame_size0_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_frame_size0_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_frame_size0_w;
wire hdmi2usbsoc_csrbank1_dma_slot0_status0_re;
wire [1:0] hdmi2usbsoc_csrbank1_dma_slot0_status0_r;
wire [1:0] hdmi2usbsoc_csrbank1_dma_slot0_status0_w;
wire hdmi2usbsoc_csrbank1_dma_slot0_address3_re;
wire [2:0] hdmi2usbsoc_csrbank1_dma_slot0_address3_r;
wire [2:0] hdmi2usbsoc_csrbank1_dma_slot0_address3_w;
wire hdmi2usbsoc_csrbank1_dma_slot0_address2_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot0_address2_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot0_address2_w;
wire hdmi2usbsoc_csrbank1_dma_slot0_address1_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot0_address1_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot0_address1_w;
wire hdmi2usbsoc_csrbank1_dma_slot0_address0_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot0_address0_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot0_address0_w;
wire hdmi2usbsoc_csrbank1_dma_slot1_status0_re;
wire [1:0] hdmi2usbsoc_csrbank1_dma_slot1_status0_r;
wire [1:0] hdmi2usbsoc_csrbank1_dma_slot1_status0_w;
wire hdmi2usbsoc_csrbank1_dma_slot1_address3_re;
wire [2:0] hdmi2usbsoc_csrbank1_dma_slot1_address3_r;
wire [2:0] hdmi2usbsoc_csrbank1_dma_slot1_address3_w;
wire hdmi2usbsoc_csrbank1_dma_slot1_address2_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot1_address2_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot1_address2_w;
wire hdmi2usbsoc_csrbank1_dma_slot1_address1_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot1_address1_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot1_address1_w;
wire hdmi2usbsoc_csrbank1_dma_slot1_address0_re;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot1_address0_r;
wire [7:0] hdmi2usbsoc_csrbank1_dma_slot1_address0_w;
wire hdmi2usbsoc_csrbank1_dma_ev_enable0_re;
wire [1:0] hdmi2usbsoc_csrbank1_dma_ev_enable0_r;
wire [1:0] hdmi2usbsoc_csrbank1_dma_ev_enable0_w;
wire hdmi2usbsoc_csrbank1_sel;
wire [13:0] hdmi2usbsoc_interface1_sram_bus_adr;
wire hdmi2usbsoc_interface1_sram_bus_we;
wire [7:0] hdmi2usbsoc_interface1_sram_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface1_sram_bus_dat_r = 8'd0;
wire [6:0] hdmi2usbsoc_sram1_adr;
wire [7:0] hdmi2usbsoc_sram1_dat_r;
wire hdmi2usbsoc_sram1_we;
wire [7:0] hdmi2usbsoc_sram1_dat_w;
wire hdmi2usbsoc_sram1_sel;
reg hdmi2usbsoc_sram1_sel_r = 1'd0;
wire [13:0] hdmi2usbsoc_interface2_bank_bus_adr;
wire hdmi2usbsoc_interface2_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface2_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface2_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank2_edid_hpd_notif_re;
wire hdmi2usbsoc_csrbank2_edid_hpd_notif_r;
wire hdmi2usbsoc_csrbank2_edid_hpd_notif_w;
wire hdmi2usbsoc_csrbank2_edid_hpd_en0_re;
wire hdmi2usbsoc_csrbank2_edid_hpd_en0_r;
wire hdmi2usbsoc_csrbank2_edid_hpd_en0_w;
wire hdmi2usbsoc_csrbank2_clocking_pll_reset0_re;
wire hdmi2usbsoc_csrbank2_clocking_pll_reset0_r;
wire hdmi2usbsoc_csrbank2_clocking_pll_reset0_w;
wire hdmi2usbsoc_csrbank2_clocking_locked_re;
wire hdmi2usbsoc_csrbank2_clocking_locked_r;
wire hdmi2usbsoc_csrbank2_clocking_locked_w;
wire hdmi2usbsoc_csrbank2_clocking_pll_adr0_re;
wire [4:0] hdmi2usbsoc_csrbank2_clocking_pll_adr0_r;
wire [4:0] hdmi2usbsoc_csrbank2_clocking_pll_adr0_w;
wire hdmi2usbsoc_csrbank2_clocking_pll_dat_r1_re;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_r1_r;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_r1_w;
wire hdmi2usbsoc_csrbank2_clocking_pll_dat_r0_re;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_r0_r;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_r0_w;
wire hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_re;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_r;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_w;
wire hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_re;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_r;
wire [7:0] hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_w;
wire hdmi2usbsoc_csrbank2_clocking_pll_drdy_re;
wire hdmi2usbsoc_csrbank2_clocking_pll_drdy_r;
wire hdmi2usbsoc_csrbank2_clocking_pll_drdy_w;
wire hdmi2usbsoc_csrbank2_data0_cap_dly_busy_re;
wire [1:0] hdmi2usbsoc_csrbank2_data0_cap_dly_busy_r;
wire [1:0] hdmi2usbsoc_csrbank2_data0_cap_dly_busy_w;
wire hdmi2usbsoc_csrbank2_data0_cap_phase_re;
wire [1:0] hdmi2usbsoc_csrbank2_data0_cap_phase_r;
wire [1:0] hdmi2usbsoc_csrbank2_data0_cap_phase_w;
wire hdmi2usbsoc_csrbank2_data0_charsync_char_synced_re;
wire hdmi2usbsoc_csrbank2_data0_charsync_char_synced_r;
wire hdmi2usbsoc_csrbank2_data0_charsync_char_synced_w;
wire hdmi2usbsoc_csrbank2_data0_charsync_ctl_pos_re;
wire [3:0] hdmi2usbsoc_csrbank2_data0_charsync_ctl_pos_r;
wire [3:0] hdmi2usbsoc_csrbank2_data0_charsync_ctl_pos_w;
wire hdmi2usbsoc_csrbank2_data0_wer_value2_re;
wire [7:0] hdmi2usbsoc_csrbank2_data0_wer_value2_r;
wire [7:0] hdmi2usbsoc_csrbank2_data0_wer_value2_w;
wire hdmi2usbsoc_csrbank2_data0_wer_value1_re;
wire [7:0] hdmi2usbsoc_csrbank2_data0_wer_value1_r;
wire [7:0] hdmi2usbsoc_csrbank2_data0_wer_value1_w;
wire hdmi2usbsoc_csrbank2_data0_wer_value0_re;
wire [7:0] hdmi2usbsoc_csrbank2_data0_wer_value0_r;
wire [7:0] hdmi2usbsoc_csrbank2_data0_wer_value0_w;
wire hdmi2usbsoc_csrbank2_data1_cap_dly_busy_re;
wire [1:0] hdmi2usbsoc_csrbank2_data1_cap_dly_busy_r;
wire [1:0] hdmi2usbsoc_csrbank2_data1_cap_dly_busy_w;
wire hdmi2usbsoc_csrbank2_data1_cap_phase_re;
wire [1:0] hdmi2usbsoc_csrbank2_data1_cap_phase_r;
wire [1:0] hdmi2usbsoc_csrbank2_data1_cap_phase_w;
wire hdmi2usbsoc_csrbank2_data1_charsync_char_synced_re;
wire hdmi2usbsoc_csrbank2_data1_charsync_char_synced_r;
wire hdmi2usbsoc_csrbank2_data1_charsync_char_synced_w;
wire hdmi2usbsoc_csrbank2_data1_charsync_ctl_pos_re;
wire [3:0] hdmi2usbsoc_csrbank2_data1_charsync_ctl_pos_r;
wire [3:0] hdmi2usbsoc_csrbank2_data1_charsync_ctl_pos_w;
wire hdmi2usbsoc_csrbank2_data1_wer_value2_re;
wire [7:0] hdmi2usbsoc_csrbank2_data1_wer_value2_r;
wire [7:0] hdmi2usbsoc_csrbank2_data1_wer_value2_w;
wire hdmi2usbsoc_csrbank2_data1_wer_value1_re;
wire [7:0] hdmi2usbsoc_csrbank2_data1_wer_value1_r;
wire [7:0] hdmi2usbsoc_csrbank2_data1_wer_value1_w;
wire hdmi2usbsoc_csrbank2_data1_wer_value0_re;
wire [7:0] hdmi2usbsoc_csrbank2_data1_wer_value0_r;
wire [7:0] hdmi2usbsoc_csrbank2_data1_wer_value0_w;
wire hdmi2usbsoc_csrbank2_data2_cap_dly_busy_re;
wire [1:0] hdmi2usbsoc_csrbank2_data2_cap_dly_busy_r;
wire [1:0] hdmi2usbsoc_csrbank2_data2_cap_dly_busy_w;
wire hdmi2usbsoc_csrbank2_data2_cap_phase_re;
wire [1:0] hdmi2usbsoc_csrbank2_data2_cap_phase_r;
wire [1:0] hdmi2usbsoc_csrbank2_data2_cap_phase_w;
wire hdmi2usbsoc_csrbank2_data2_charsync_char_synced_re;
wire hdmi2usbsoc_csrbank2_data2_charsync_char_synced_r;
wire hdmi2usbsoc_csrbank2_data2_charsync_char_synced_w;
wire hdmi2usbsoc_csrbank2_data2_charsync_ctl_pos_re;
wire [3:0] hdmi2usbsoc_csrbank2_data2_charsync_ctl_pos_r;
wire [3:0] hdmi2usbsoc_csrbank2_data2_charsync_ctl_pos_w;
wire hdmi2usbsoc_csrbank2_data2_wer_value2_re;
wire [7:0] hdmi2usbsoc_csrbank2_data2_wer_value2_r;
wire [7:0] hdmi2usbsoc_csrbank2_data2_wer_value2_w;
wire hdmi2usbsoc_csrbank2_data2_wer_value1_re;
wire [7:0] hdmi2usbsoc_csrbank2_data2_wer_value1_r;
wire [7:0] hdmi2usbsoc_csrbank2_data2_wer_value1_w;
wire hdmi2usbsoc_csrbank2_data2_wer_value0_re;
wire [7:0] hdmi2usbsoc_csrbank2_data2_wer_value0_r;
wire [7:0] hdmi2usbsoc_csrbank2_data2_wer_value0_w;
wire hdmi2usbsoc_csrbank2_chansync_channels_synced_re;
wire hdmi2usbsoc_csrbank2_chansync_channels_synced_r;
wire hdmi2usbsoc_csrbank2_chansync_channels_synced_w;
wire hdmi2usbsoc_csrbank2_resdetection_hres1_re;
wire [2:0] hdmi2usbsoc_csrbank2_resdetection_hres1_r;
wire [2:0] hdmi2usbsoc_csrbank2_resdetection_hres1_w;
wire hdmi2usbsoc_csrbank2_resdetection_hres0_re;
wire [7:0] hdmi2usbsoc_csrbank2_resdetection_hres0_r;
wire [7:0] hdmi2usbsoc_csrbank2_resdetection_hres0_w;
wire hdmi2usbsoc_csrbank2_resdetection_vres1_re;
wire [2:0] hdmi2usbsoc_csrbank2_resdetection_vres1_r;
wire [2:0] hdmi2usbsoc_csrbank2_resdetection_vres1_w;
wire hdmi2usbsoc_csrbank2_resdetection_vres0_re;
wire [7:0] hdmi2usbsoc_csrbank2_resdetection_vres0_r;
wire [7:0] hdmi2usbsoc_csrbank2_resdetection_vres0_w;
wire hdmi2usbsoc_csrbank2_dma_frame_size3_re;
wire [2:0] hdmi2usbsoc_csrbank2_dma_frame_size3_r;
wire [2:0] hdmi2usbsoc_csrbank2_dma_frame_size3_w;
wire hdmi2usbsoc_csrbank2_dma_frame_size2_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_frame_size2_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_frame_size2_w;
wire hdmi2usbsoc_csrbank2_dma_frame_size1_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_frame_size1_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_frame_size1_w;
wire hdmi2usbsoc_csrbank2_dma_frame_size0_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_frame_size0_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_frame_size0_w;
wire hdmi2usbsoc_csrbank2_dma_slot0_status0_re;
wire [1:0] hdmi2usbsoc_csrbank2_dma_slot0_status0_r;
wire [1:0] hdmi2usbsoc_csrbank2_dma_slot0_status0_w;
wire hdmi2usbsoc_csrbank2_dma_slot0_address3_re;
wire [2:0] hdmi2usbsoc_csrbank2_dma_slot0_address3_r;
wire [2:0] hdmi2usbsoc_csrbank2_dma_slot0_address3_w;
wire hdmi2usbsoc_csrbank2_dma_slot0_address2_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot0_address2_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot0_address2_w;
wire hdmi2usbsoc_csrbank2_dma_slot0_address1_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot0_address1_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot0_address1_w;
wire hdmi2usbsoc_csrbank2_dma_slot0_address0_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot0_address0_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot0_address0_w;
wire hdmi2usbsoc_csrbank2_dma_slot1_status0_re;
wire [1:0] hdmi2usbsoc_csrbank2_dma_slot1_status0_r;
wire [1:0] hdmi2usbsoc_csrbank2_dma_slot1_status0_w;
wire hdmi2usbsoc_csrbank2_dma_slot1_address3_re;
wire [2:0] hdmi2usbsoc_csrbank2_dma_slot1_address3_r;
wire [2:0] hdmi2usbsoc_csrbank2_dma_slot1_address3_w;
wire hdmi2usbsoc_csrbank2_dma_slot1_address2_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot1_address2_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot1_address2_w;
wire hdmi2usbsoc_csrbank2_dma_slot1_address1_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot1_address1_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot1_address1_w;
wire hdmi2usbsoc_csrbank2_dma_slot1_address0_re;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot1_address0_r;
wire [7:0] hdmi2usbsoc_csrbank2_dma_slot1_address0_w;
wire hdmi2usbsoc_csrbank2_dma_ev_enable0_re;
wire [1:0] hdmi2usbsoc_csrbank2_dma_ev_enable0_r;
wire [1:0] hdmi2usbsoc_csrbank2_dma_ev_enable0_w;
wire hdmi2usbsoc_csrbank2_sel;
wire [13:0] hdmi2usbsoc_interface3_bank_bus_adr;
wire hdmi2usbsoc_interface3_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface3_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface3_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank3_core_underflow_enable0_re;
wire hdmi2usbsoc_csrbank3_core_underflow_enable0_r;
wire hdmi2usbsoc_csrbank3_core_underflow_enable0_w;
wire hdmi2usbsoc_csrbank3_core_underflow_counter3_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter3_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter3_w;
wire hdmi2usbsoc_csrbank3_core_underflow_counter2_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter2_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter2_w;
wire hdmi2usbsoc_csrbank3_core_underflow_counter1_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter1_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter1_w;
wire hdmi2usbsoc_csrbank3_core_underflow_counter0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_underflow_counter0_w;
wire hdmi2usbsoc_csrbank3_core_initiator_enable0_re;
wire hdmi2usbsoc_csrbank3_core_initiator_enable0_r;
wire hdmi2usbsoc_csrbank3_core_initiator_enable0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_hres_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_hres1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hres1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hres1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_hres0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hres0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hres0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_start_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_end_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_hscan_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_hscan1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hscan1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_hscan1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_hscan0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hscan0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_hscan0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_vres_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_vres1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vres1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vres1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_vres0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vres0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vres0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_start_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_end_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_w;
reg [3:0] hdmi2usbsoc_csrbank3_core_initiator_vscan_backstore = 4'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_vscan1_re;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vscan1_r;
wire [3:0] hdmi2usbsoc_csrbank3_core_initiator_vscan1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_vscan0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vscan0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_vscan0_w;
reg [23:0] hdmi2usbsoc_csrbank3_core_initiator_base_backstore = 24'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_base3_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base3_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base3_w;
wire hdmi2usbsoc_csrbank3_core_initiator_base2_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base2_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base2_w;
wire hdmi2usbsoc_csrbank3_core_initiator_base1_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base1_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_base0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_base0_w;
reg [23:0] hdmi2usbsoc_csrbank3_core_initiator_length_backstore = 24'd0;
wire hdmi2usbsoc_csrbank3_core_initiator_length3_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length3_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length3_w;
wire hdmi2usbsoc_csrbank3_core_initiator_length2_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length2_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length2_w;
wire hdmi2usbsoc_csrbank3_core_initiator_length1_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length1_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length1_w;
wire hdmi2usbsoc_csrbank3_core_initiator_length0_re;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length0_r;
wire [7:0] hdmi2usbsoc_csrbank3_core_initiator_length0_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_re;
wire [1:0] hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_r;
wire [1:0] hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_re;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_r;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_status_re;
wire [3:0] hdmi2usbsoc_csrbank3_driver_clocking_status_r;
wire [3:0] hdmi2usbsoc_csrbank3_driver_clocking_status_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_re;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_r;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_re;
wire [4:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_r;
wire [4:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r1_re;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r1_r;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r1_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r0_re;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r0_r;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r0_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_re;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_r;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_re;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_r;
wire [7:0] hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_w;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_drdy_re;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_drdy_r;
wire hdmi2usbsoc_csrbank3_driver_clocking_pll_drdy_w;
wire hdmi2usbsoc_csrbank3_sel;
wire [13:0] hdmi2usbsoc_interface4_bank_bus_adr;
wire hdmi2usbsoc_interface4_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface4_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface4_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank4_core_underflow_enable0_re;
wire hdmi2usbsoc_csrbank4_core_underflow_enable0_r;
wire hdmi2usbsoc_csrbank4_core_underflow_enable0_w;
wire hdmi2usbsoc_csrbank4_core_underflow_counter3_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter3_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter3_w;
wire hdmi2usbsoc_csrbank4_core_underflow_counter2_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter2_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter2_w;
wire hdmi2usbsoc_csrbank4_core_underflow_counter1_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter1_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter1_w;
wire hdmi2usbsoc_csrbank4_core_underflow_counter0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_underflow_counter0_w;
wire hdmi2usbsoc_csrbank4_core_initiator_enable0_re;
wire hdmi2usbsoc_csrbank4_core_initiator_enable0_r;
wire hdmi2usbsoc_csrbank4_core_initiator_enable0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_hres_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_hres1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hres1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hres1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_hres0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hres0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hres0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_start_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_end_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_hscan_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_hscan1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hscan1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_hscan1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_hscan0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hscan0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_hscan0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_vres_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_vres1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vres1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vres1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_vres0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vres0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vres0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_start_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_end_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_w;
reg [3:0] hdmi2usbsoc_csrbank4_core_initiator_vscan_backstore = 4'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_vscan1_re;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vscan1_r;
wire [3:0] hdmi2usbsoc_csrbank4_core_initiator_vscan1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_vscan0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vscan0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_vscan0_w;
reg [23:0] hdmi2usbsoc_csrbank4_core_initiator_base_backstore = 24'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_base3_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base3_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base3_w;
wire hdmi2usbsoc_csrbank4_core_initiator_base2_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base2_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base2_w;
wire hdmi2usbsoc_csrbank4_core_initiator_base1_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base1_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_base0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_base0_w;
reg [23:0] hdmi2usbsoc_csrbank4_core_initiator_length_backstore = 24'd0;
wire hdmi2usbsoc_csrbank4_core_initiator_length3_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length3_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length3_w;
wire hdmi2usbsoc_csrbank4_core_initiator_length2_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length2_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length2_w;
wire hdmi2usbsoc_csrbank4_core_initiator_length1_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length1_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length1_w;
wire hdmi2usbsoc_csrbank4_core_initiator_length0_re;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length0_r;
wire [7:0] hdmi2usbsoc_csrbank4_core_initiator_length0_w;
wire hdmi2usbsoc_csrbank4_sel;
wire [13:0] hdmi2usbsoc_interface2_sram_bus_adr;
wire hdmi2usbsoc_interface2_sram_bus_we;
wire [7:0] hdmi2usbsoc_interface2_sram_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface2_sram_bus_dat_r = 8'd0;
wire [3:0] hdmi2usbsoc_sram2_adr;
wire [7:0] hdmi2usbsoc_sram2_dat_r;
wire hdmi2usbsoc_sram2_sel;
reg hdmi2usbsoc_sram2_sel_r = 1'd0;
wire [13:0] hdmi2usbsoc_interface5_bank_bus_adr;
wire hdmi2usbsoc_interface5_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface5_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface5_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank5_dna_id7_re;
wire hdmi2usbsoc_csrbank5_dna_id7_r;
wire hdmi2usbsoc_csrbank5_dna_id7_w;
wire hdmi2usbsoc_csrbank5_dna_id6_re;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id6_r;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id6_w;
wire hdmi2usbsoc_csrbank5_dna_id5_re;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id5_r;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id5_w;
wire hdmi2usbsoc_csrbank5_dna_id4_re;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id4_r;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id4_w;
wire hdmi2usbsoc_csrbank5_dna_id3_re;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id3_r;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id3_w;
wire hdmi2usbsoc_csrbank5_dna_id2_re;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id2_r;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id2_w;
wire hdmi2usbsoc_csrbank5_dna_id1_re;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id1_r;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id1_w;
wire hdmi2usbsoc_csrbank5_dna_id0_re;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id0_r;
wire [7:0] hdmi2usbsoc_csrbank5_dna_id0_w;
wire hdmi2usbsoc_csrbank5_git_commit19_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit19_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit19_w;
wire hdmi2usbsoc_csrbank5_git_commit18_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit18_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit18_w;
wire hdmi2usbsoc_csrbank5_git_commit17_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit17_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit17_w;
wire hdmi2usbsoc_csrbank5_git_commit16_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit16_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit16_w;
wire hdmi2usbsoc_csrbank5_git_commit15_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit15_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit15_w;
wire hdmi2usbsoc_csrbank5_git_commit14_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit14_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit14_w;
wire hdmi2usbsoc_csrbank5_git_commit13_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit13_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit13_w;
wire hdmi2usbsoc_csrbank5_git_commit12_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit12_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit12_w;
wire hdmi2usbsoc_csrbank5_git_commit11_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit11_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit11_w;
wire hdmi2usbsoc_csrbank5_git_commit10_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit10_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit10_w;
wire hdmi2usbsoc_csrbank5_git_commit9_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit9_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit9_w;
wire hdmi2usbsoc_csrbank5_git_commit8_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit8_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit8_w;
wire hdmi2usbsoc_csrbank5_git_commit7_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit7_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit7_w;
wire hdmi2usbsoc_csrbank5_git_commit6_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit6_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit6_w;
wire hdmi2usbsoc_csrbank5_git_commit5_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit5_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit5_w;
wire hdmi2usbsoc_csrbank5_git_commit4_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit4_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit4_w;
wire hdmi2usbsoc_csrbank5_git_commit3_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit3_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit3_w;
wire hdmi2usbsoc_csrbank5_git_commit2_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit2_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit2_w;
wire hdmi2usbsoc_csrbank5_git_commit1_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit1_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit1_w;
wire hdmi2usbsoc_csrbank5_git_commit0_re;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit0_r;
wire [7:0] hdmi2usbsoc_csrbank5_git_commit0_w;
wire hdmi2usbsoc_csrbank5_platform_platform7_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform7_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform7_w;
wire hdmi2usbsoc_csrbank5_platform_platform6_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform6_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform6_w;
wire hdmi2usbsoc_csrbank5_platform_platform5_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform5_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform5_w;
wire hdmi2usbsoc_csrbank5_platform_platform4_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform4_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform4_w;
wire hdmi2usbsoc_csrbank5_platform_platform3_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform3_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform3_w;
wire hdmi2usbsoc_csrbank5_platform_platform2_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform2_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform2_w;
wire hdmi2usbsoc_csrbank5_platform_platform1_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform1_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform1_w;
wire hdmi2usbsoc_csrbank5_platform_platform0_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform0_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_platform0_w;
wire hdmi2usbsoc_csrbank5_platform_target7_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target7_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target7_w;
wire hdmi2usbsoc_csrbank5_platform_target6_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target6_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target6_w;
wire hdmi2usbsoc_csrbank5_platform_target5_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target5_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target5_w;
wire hdmi2usbsoc_csrbank5_platform_target4_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target4_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target4_w;
wire hdmi2usbsoc_csrbank5_platform_target3_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target3_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target3_w;
wire hdmi2usbsoc_csrbank5_platform_target2_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target2_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target2_w;
wire hdmi2usbsoc_csrbank5_platform_target1_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target1_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target1_w;
wire hdmi2usbsoc_csrbank5_platform_target0_re;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target0_r;
wire [7:0] hdmi2usbsoc_csrbank5_platform_target0_w;
wire hdmi2usbsoc_csrbank5_sel;
wire [13:0] hdmi2usbsoc_interface6_bank_bus_adr;
wire hdmi2usbsoc_interface6_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface6_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface6_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank6_dfii_control0_re;
wire [3:0] hdmi2usbsoc_csrbank6_dfii_control0_r;
wire [3:0] hdmi2usbsoc_csrbank6_dfii_control0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_command0_re;
wire [5:0] hdmi2usbsoc_csrbank6_dfii_pi0_command0_r;
wire [5:0] hdmi2usbsoc_csrbank6_dfii_pi0_command0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_address1_re;
wire [4:0] hdmi2usbsoc_csrbank6_dfii_pi0_address1_r;
wire [4:0] hdmi2usbsoc_csrbank6_dfii_pi0_address1_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_address0_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_address0_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_address0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_re;
wire [2:0] hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_r;
wire [2:0] hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_rddata3_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata3_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata3_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_rddata2_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata2_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata2_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_rddata1_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata1_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata1_w;
wire hdmi2usbsoc_csrbank6_dfii_pi0_rddata0_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata0_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi0_rddata0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_command0_re;
wire [5:0] hdmi2usbsoc_csrbank6_dfii_pi1_command0_r;
wire [5:0] hdmi2usbsoc_csrbank6_dfii_pi1_command0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_address1_re;
wire [4:0] hdmi2usbsoc_csrbank6_dfii_pi1_address1_r;
wire [4:0] hdmi2usbsoc_csrbank6_dfii_pi1_address1_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_address0_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_address0_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_address0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_re;
wire [2:0] hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_r;
wire [2:0] hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_rddata3_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata3_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata3_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_rddata2_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata2_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata2_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_rddata1_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata1_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata1_w;
wire hdmi2usbsoc_csrbank6_dfii_pi1_rddata0_re;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata0_r;
wire [7:0] hdmi2usbsoc_csrbank6_dfii_pi1_rddata0_w;
wire hdmi2usbsoc_csrbank6_controller_bandwidth_nreads2_re;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nreads2_r;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nreads2_w;
wire hdmi2usbsoc_csrbank6_controller_bandwidth_nreads1_re;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nreads1_r;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nreads1_w;
wire hdmi2usbsoc_csrbank6_controller_bandwidth_nreads0_re;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nreads0_r;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nreads0_w;
wire hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites2_re;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites2_r;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites2_w;
wire hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites1_re;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites1_r;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites1_w;
wire hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites0_re;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites0_r;
wire [7:0] hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites0_w;
wire hdmi2usbsoc_csrbank6_controller_bandwidth_data_width_re;
wire [6:0] hdmi2usbsoc_csrbank6_controller_bandwidth_data_width_r;
wire [6:0] hdmi2usbsoc_csrbank6_controller_bandwidth_data_width_w;
wire hdmi2usbsoc_csrbank6_sel;
wire [13:0] hdmi2usbsoc_interface7_bank_bus_adr;
wire hdmi2usbsoc_interface7_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface7_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface7_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank7_bitbang0_re;
wire [3:0] hdmi2usbsoc_csrbank7_bitbang0_r;
wire [3:0] hdmi2usbsoc_csrbank7_bitbang0_w;
wire hdmi2usbsoc_csrbank7_miso_re;
wire hdmi2usbsoc_csrbank7_miso_r;
wire hdmi2usbsoc_csrbank7_miso_w;
wire hdmi2usbsoc_csrbank7_bitbang_en0_re;
wire hdmi2usbsoc_csrbank7_bitbang_en0_r;
wire hdmi2usbsoc_csrbank7_bitbang_en0_w;
wire hdmi2usbsoc_csrbank7_sel;
wire [13:0] hdmi2usbsoc_interface8_bank_bus_adr;
wire hdmi2usbsoc_interface8_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface8_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface8_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank8_load3_re;
wire [7:0] hdmi2usbsoc_csrbank8_load3_r;
wire [7:0] hdmi2usbsoc_csrbank8_load3_w;
wire hdmi2usbsoc_csrbank8_load2_re;
wire [7:0] hdmi2usbsoc_csrbank8_load2_r;
wire [7:0] hdmi2usbsoc_csrbank8_load2_w;
wire hdmi2usbsoc_csrbank8_load1_re;
wire [7:0] hdmi2usbsoc_csrbank8_load1_r;
wire [7:0] hdmi2usbsoc_csrbank8_load1_w;
wire hdmi2usbsoc_csrbank8_load0_re;
wire [7:0] hdmi2usbsoc_csrbank8_load0_r;
wire [7:0] hdmi2usbsoc_csrbank8_load0_w;
wire hdmi2usbsoc_csrbank8_reload3_re;
wire [7:0] hdmi2usbsoc_csrbank8_reload3_r;
wire [7:0] hdmi2usbsoc_csrbank8_reload3_w;
wire hdmi2usbsoc_csrbank8_reload2_re;
wire [7:0] hdmi2usbsoc_csrbank8_reload2_r;
wire [7:0] hdmi2usbsoc_csrbank8_reload2_w;
wire hdmi2usbsoc_csrbank8_reload1_re;
wire [7:0] hdmi2usbsoc_csrbank8_reload1_r;
wire [7:0] hdmi2usbsoc_csrbank8_reload1_w;
wire hdmi2usbsoc_csrbank8_reload0_re;
wire [7:0] hdmi2usbsoc_csrbank8_reload0_r;
wire [7:0] hdmi2usbsoc_csrbank8_reload0_w;
wire hdmi2usbsoc_csrbank8_en0_re;
wire hdmi2usbsoc_csrbank8_en0_r;
wire hdmi2usbsoc_csrbank8_en0_w;
wire hdmi2usbsoc_csrbank8_value3_re;
wire [7:0] hdmi2usbsoc_csrbank8_value3_r;
wire [7:0] hdmi2usbsoc_csrbank8_value3_w;
wire hdmi2usbsoc_csrbank8_value2_re;
wire [7:0] hdmi2usbsoc_csrbank8_value2_r;
wire [7:0] hdmi2usbsoc_csrbank8_value2_w;
wire hdmi2usbsoc_csrbank8_value1_re;
wire [7:0] hdmi2usbsoc_csrbank8_value1_r;
wire [7:0] hdmi2usbsoc_csrbank8_value1_w;
wire hdmi2usbsoc_csrbank8_value0_re;
wire [7:0] hdmi2usbsoc_csrbank8_value0_r;
wire [7:0] hdmi2usbsoc_csrbank8_value0_w;
wire hdmi2usbsoc_csrbank8_ev_enable0_re;
wire hdmi2usbsoc_csrbank8_ev_enable0_r;
wire hdmi2usbsoc_csrbank8_ev_enable0_w;
wire hdmi2usbsoc_csrbank8_sel;
wire [13:0] hdmi2usbsoc_interface9_bank_bus_adr;
wire hdmi2usbsoc_interface9_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface9_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface9_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank9_txfull_re;
wire hdmi2usbsoc_csrbank9_txfull_r;
wire hdmi2usbsoc_csrbank9_txfull_w;
wire hdmi2usbsoc_csrbank9_rxempty_re;
wire hdmi2usbsoc_csrbank9_rxempty_r;
wire hdmi2usbsoc_csrbank9_rxempty_w;
wire hdmi2usbsoc_csrbank9_ev_enable0_re;
wire [1:0] hdmi2usbsoc_csrbank9_ev_enable0_r;
wire [1:0] hdmi2usbsoc_csrbank9_ev_enable0_w;
wire hdmi2usbsoc_csrbank9_sel;
wire [13:0] hdmi2usbsoc_interface10_bank_bus_adr;
wire hdmi2usbsoc_interface10_bank_bus_we;
wire [7:0] hdmi2usbsoc_interface10_bank_bus_dat_w;
reg [7:0] hdmi2usbsoc_interface10_bank_bus_dat_r = 8'd0;
wire hdmi2usbsoc_csrbank10_tuning_word3_re;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word3_r;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word3_w;
wire hdmi2usbsoc_csrbank10_tuning_word2_re;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word2_r;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word2_w;
wire hdmi2usbsoc_csrbank10_tuning_word1_re;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word1_r;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word1_w;
wire hdmi2usbsoc_csrbank10_tuning_word0_re;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word0_r;
wire [7:0] hdmi2usbsoc_csrbank10_tuning_word0_w;
wire hdmi2usbsoc_csrbank10_sel;
wire [15:0] slice_proxy0;
wire [15:0] slice_proxy1;
wire [15:0] slice_proxy2;
wire [15:0] slice_proxy3;
wire [15:0] slice_proxy4;
wire [15:0] slice_proxy5;
wire [15:0] slice_proxy6;
wire [15:0] slice_proxy7;
wire [15:0] slice_proxy8;
wire [15:0] slice_proxy9;
wire [15:0] slice_proxy10;
wire [15:0] slice_proxy11;
wire [15:0] slice_proxy12;
wire [15:0] slice_proxy13;
wire [15:0] slice_proxy14;
wire [15:0] slice_proxy15;
wire [15:0] slice_proxy16;
wire [15:0] slice_proxy17;
wire [15:0] slice_proxy18;
wire [15:0] slice_proxy19;
wire [15:0] slice_proxy20;
wire [15:0] slice_proxy21;
wire [15:0] slice_proxy22;
wire [15:0] slice_proxy23;
wire [15:0] slice_proxy24;
wire [15:0] slice_proxy25;
wire [15:0] slice_proxy26;
wire [15:0] slice_proxy27;
wire [15:0] slice_proxy28;
wire [15:0] slice_proxy29;
wire [15:0] slice_proxy30;
wire [15:0] slice_proxy31;
wire [15:0] slice_proxy32;
wire [15:0] slice_proxy33;
wire [15:0] slice_proxy34;
wire [15:0] slice_proxy35;
wire [15:0] slice_proxy36;
wire [15:0] slice_proxy37;
wire [15:0] slice_proxy38;
wire [15:0] slice_proxy39;
wire [15:0] slice_proxy40;
wire [15:0] slice_proxy41;
wire [15:0] slice_proxy42;
wire [15:0] slice_proxy43;
wire [15:0] slice_proxy44;
wire [15:0] slice_proxy45;
wire [15:0] slice_proxy46;
wire [15:0] slice_proxy47;
wire [15:0] slice_proxy48;
wire [15:0] slice_proxy49;
wire [15:0] slice_proxy50;
wire [15:0] slice_proxy51;
wire [15:0] slice_proxy52;
wire [15:0] slice_proxy53;
wire [15:0] slice_proxy54;
wire [15:0] slice_proxy55;
wire [15:0] slice_proxy56;
wire [15:0] slice_proxy57;
wire [15:0] slice_proxy58;
wire [15:0] slice_proxy59;
wire [15:0] slice_proxy60;
wire [15:0] slice_proxy61;
wire [15:0] slice_proxy62;
wire [15:0] slice_proxy63;
wire [1:0] slice_proxy64;
wire [1:0] slice_proxy65;
wire [1:0] slice_proxy66;
wire [1:0] slice_proxy67;
wire [1:0] slice_proxy68;
wire [1:0] slice_proxy69;
wire [1:0] slice_proxy70;
wire [1:0] slice_proxy71;
reg comb_rhs_array_muxed0 = 1'd0;
reg [12:0] comb_rhs_array_muxed1 = 13'd0;
reg [2:0] comb_rhs_array_muxed2 = 3'd0;
reg comb_rhs_array_muxed3 = 1'd0;
reg comb_rhs_array_muxed4 = 1'd0;
reg comb_rhs_array_muxed5 = 1'd0;
reg comb_t_array_muxed0 = 1'd0;
reg comb_t_array_muxed1 = 1'd0;
reg comb_t_array_muxed2 = 1'd0;
reg comb_rhs_array_muxed6 = 1'd0;
reg [12:0] comb_rhs_array_muxed7 = 13'd0;
reg [2:0] comb_rhs_array_muxed8 = 3'd0;
reg comb_rhs_array_muxed9 = 1'd0;
reg comb_rhs_array_muxed10 = 1'd0;
reg comb_rhs_array_muxed11 = 1'd0;
reg comb_t_array_muxed3 = 1'd0;
reg comb_t_array_muxed4 = 1'd0;
reg comb_t_array_muxed5 = 1'd0;
reg [20:0] comb_rhs_array_muxed12 = 21'd0;
reg comb_rhs_array_muxed13 = 1'd0;
reg comb_rhs_array_muxed14 = 1'd0;
reg [20:0] comb_rhs_array_muxed15 = 21'd0;
reg comb_rhs_array_muxed16 = 1'd0;
reg comb_rhs_array_muxed17 = 1'd0;
reg [20:0] comb_rhs_array_muxed18 = 21'd0;
reg comb_rhs_array_muxed19 = 1'd0;
reg comb_rhs_array_muxed20 = 1'd0;
reg [20:0] comb_rhs_array_muxed21 = 21'd0;
reg comb_rhs_array_muxed22 = 1'd0;
reg comb_rhs_array_muxed23 = 1'd0;
reg [20:0] comb_rhs_array_muxed24 = 21'd0;
reg comb_rhs_array_muxed25 = 1'd0;
reg comb_rhs_array_muxed26 = 1'd0;
reg [20:0] comb_rhs_array_muxed27 = 21'd0;
reg comb_rhs_array_muxed28 = 1'd0;
reg comb_rhs_array_muxed29 = 1'd0;
reg [20:0] comb_rhs_array_muxed30 = 21'd0;
reg comb_rhs_array_muxed31 = 1'd0;
reg comb_rhs_array_muxed32 = 1'd0;
reg [20:0] comb_rhs_array_muxed33 = 21'd0;
reg comb_rhs_array_muxed34 = 1'd0;
reg comb_rhs_array_muxed35 = 1'd0;
reg [23:0] comb_rhs_array_muxed36 = 24'd0;
reg comb_rhs_array_muxed37 = 1'd0;
reg [23:0] comb_rhs_array_muxed38 = 24'd0;
reg comb_rhs_array_muxed39 = 1'd0;
reg [29:0] comb_rhs_array_muxed40 = 30'd0;
reg [31:0] comb_rhs_array_muxed41 = 32'd0;
reg [3:0] comb_rhs_array_muxed42 = 4'd0;
reg comb_rhs_array_muxed43 = 1'd0;
reg comb_rhs_array_muxed44 = 1'd0;
reg comb_rhs_array_muxed45 = 1'd0;
reg [2:0] comb_rhs_array_muxed46 = 3'd0;
reg [1:0] comb_rhs_array_muxed47 = 2'd0;
reg [29:0] comb_rhs_array_muxed48 = 30'd0;
reg [31:0] comb_rhs_array_muxed49 = 32'd0;
reg [3:0] comb_rhs_array_muxed50 = 4'd0;
reg comb_rhs_array_muxed51 = 1'd0;
reg comb_rhs_array_muxed52 = 1'd0;
reg comb_rhs_array_muxed53 = 1'd0;
reg [2:0] comb_rhs_array_muxed54 = 3'd0;
reg [1:0] comb_rhs_array_muxed55 = 2'd0;
reg [9:0] sync_f_array_muxed0 = 10'd0;
reg [9:0] sync_f_array_muxed1 = 10'd0;
reg [9:0] sync_f_array_muxed2 = 10'd0;
reg [9:0] sync_f_array_muxed3 = 10'd0;
reg [9:0] sync_f_array_muxed4 = 10'd0;
reg [9:0] sync_f_array_muxed5 = 10'd0;
reg [12:0] sync_rhs_array_muxed0 = 13'd0;
reg [2:0] sync_rhs_array_muxed1 = 3'd0;
reg sync_rhs_array_muxed2 = 1'd0;
reg sync_rhs_array_muxed3 = 1'd0;
reg sync_rhs_array_muxed4 = 1'd0;
reg sync_rhs_array_muxed5 = 1'd0;
reg sync_rhs_array_muxed6 = 1'd0;
reg [12:0] sync_rhs_array_muxed7 = 13'd0;
reg [2:0] sync_rhs_array_muxed8 = 3'd0;
reg sync_rhs_array_muxed9 = 1'd0;
reg sync_rhs_array_muxed10 = 1'd0;
reg sync_rhs_array_muxed11 = 1'd0;
reg sync_rhs_array_muxed12 = 1'd0;
reg sync_rhs_array_muxed13 = 1'd0;
reg [12:0] sync_rhs_array_muxed14 = 13'd0;
reg [2:0] sync_rhs_array_muxed15 = 3'd0;
reg sync_rhs_array_muxed16 = 1'd0;
reg sync_rhs_array_muxed17 = 1'd0;
reg sync_rhs_array_muxed18 = 1'd0;
reg sync_rhs_array_muxed19 = 1'd0;
reg sync_rhs_array_muxed20 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl0_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl0_regs1 = 1'd0;
wire xilinxasyncresetsynchronizerimpl0;
wire xilinxasyncresetsynchronizerimpl0_rst_meta;
wire xilinxasyncresetsynchronizerimpl1;
wire xilinxasyncresetsynchronizerimpl1_rst_meta;
wire xilinxasyncresetsynchronizerimpl2;
wire xilinxasyncresetsynchronizerimpl2_rst_meta;
wire xilinxasyncresetsynchronizerimpl3_rst_meta;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl1_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl1_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl2_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl2_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl3_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl3_regs1 = 1'd0;
wire xilinxasyncresetsynchronizerimpl4;
wire xilinxasyncresetsynchronizerimpl4_rst_meta;
wire xilinxasyncresetsynchronizerimpl5;
wire xilinxasyncresetsynchronizerimpl5_rst_meta;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl4_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl4_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl5_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl5_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl6_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl6_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl7_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl7_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl8_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl8_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl9_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl9_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl10_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl10_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl11_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl11_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl12_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl12_regs1 = 2'd0;
wire xilinxmultiregimpl12;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl13_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl13_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl14_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl14_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl15_regs0 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl15_regs1 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl16_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl16_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl17_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl17_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl18_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl18_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl19_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl19_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl20_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl20_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl21_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl21_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl22_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl22_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl23_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl23_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl24_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl24_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl25_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl25_regs1 = 2'd0;
wire xilinxmultiregimpl25;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl26_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl26_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl27_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl27_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl28_regs0 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl28_regs1 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl29_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl29_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl30_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl30_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl31_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl31_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl32_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl32_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl33_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl33_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl34_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl34_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl35_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl35_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl36_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl36_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl37_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl37_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl38_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl38_regs1 = 2'd0;
wire xilinxmultiregimpl38;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl39_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl39_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl40_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl40_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl41_regs0 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl41_regs1 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl42_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl42_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl43_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl43_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl44_regs0 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl44_regs1 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl45_regs0 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl45_regs1 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl46_regs0 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl46_regs1 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl47_regs0 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl47_regs1 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl48_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl48_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl49_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl49_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl50_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl50_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl51_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl51_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl52_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl52_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl53_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl53_regs1 = 1'd0;
wire xilinxasyncresetsynchronizerimpl6;
wire xilinxasyncresetsynchronizerimpl6_rst_meta;
wire xilinxasyncresetsynchronizerimpl7;
wire xilinxasyncresetsynchronizerimpl7_rst_meta;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl54_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl54_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl55_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl55_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl56_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl56_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl57_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl57_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl58_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl58_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl59_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl59_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl60_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl60_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl61_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl61_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl62_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl62_regs1 = 2'd0;
wire xilinxmultiregimpl62;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl63_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl63_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl64_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl64_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl65_regs0 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl65_regs1 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl66_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl66_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl67_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl67_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl68_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl68_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl69_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl69_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl70_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl70_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl71_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl71_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl72_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl72_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl73_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl73_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl74_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl74_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl75_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl75_regs1 = 2'd0;
wire xilinxmultiregimpl75;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl76_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl76_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl77_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl77_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl78_regs0 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl78_regs1 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl79_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl79_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl80_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl80_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl81_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl81_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl82_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl82_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl83_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl83_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl84_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl84_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl85_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl85_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl86_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl86_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl87_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl87_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl88_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl88_regs1 = 2'd0;
wire xilinxmultiregimpl88;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl89_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl89_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl90_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl90_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl91_regs0 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [3:0] xilinxmultiregimpl91_regs1 = 4'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl92_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl92_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl93_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl93_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl94_regs0 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl94_regs1 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl95_regs0 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [10:0] xilinxmultiregimpl95_regs1 = 11'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl96_regs0 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl96_regs1 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl97_regs0 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [9:0] xilinxmultiregimpl97_regs1 = 10'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl98_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl98_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl99_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl99_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl100_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl100_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl101_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl101_regs1 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl102_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl102_regs1 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl103_regs0 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl103_regs1 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl104_regs0 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl104_regs1 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl105_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl105_regs1 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl106_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl106_regs1 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl107_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl107_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl108_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl108_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl109_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl109_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl110_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl110_regs1 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl111_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl111_regs1 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl112_regs0 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl112_regs1 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl113_regs0 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [4:0] xilinxmultiregimpl113_regs1 = 5'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl114_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl114_regs1 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl115_regs0 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [1:0] xilinxmultiregimpl115_regs1 = 2'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl116_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl116_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl117_regs0 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg xilinxmultiregimpl117_regs1 = 1'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl118_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl118_regs1 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl119_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl119_regs1 = 3'd0;
wire xilinxasyncresetsynchronizerimpl8_rst_meta;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl120_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl120_regs1 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl121_regs0 = 3'd0;
(* register_balancing = "no", shreg_extract = "no" *) reg [2:0] xilinxmultiregimpl121_regs1 = 3'd0;


// Adding a dummy event (using a dummy signal 'dummy_s') to get the simulator
// to run the combinatorial process once at the beginning.
// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign hdmi2usbsoc_ddrphy_clk4x_wr_strb = hdmi2usbsoc_crg_clk4x_wr_strb;
assign hdmi2usbsoc_ddrphy_clk4x_rd_strb = hdmi2usbsoc_crg_clk4x_rd_strb;
assign encoder_cdc_sink_valid = encoder_reader_source_valid;
assign encoder_reader_source_ready = encoder_cdc_sink_ready;
assign encoder_cdc_sink_first = encoder_reader_source_first;
assign encoder_cdc_sink_last = encoder_reader_source_last;
assign encoder_cdc_sink_payload_data = encoder_reader_source_payload_data;
assign encoderbuffer_sink_valid = encoder_cdc_source_valid;
assign encoder_cdc_source_ready = encoderbuffer_sink_ready;
assign encoderbuffer_sink_first = encoder_cdc_source_first;
assign encoderbuffer_sink_last = encoder_cdc_source_last;
assign encoderbuffer_sink_payload_data = encoder_cdc_source_payload_data;
assign encoder_sink_sink_valid0 = encoderbuffer_source_valid;
assign encoderbuffer_source_ready = encoder_sink_sink_ready0;
assign encoder_sink_sink_first0 = encoderbuffer_source_first;
assign encoder_sink_sink_last0 = encoderbuffer_source_last;
assign encoder_sink_sink_payload_data = encoderbuffer_source_payload_data;
assign encoder_streamer_sink_sink_valid = encoder_source_source_valid0;
assign encoder_source_source_ready0 = encoder_streamer_sink_sink_ready;
assign encoder_streamer_sink_sink_first = encoder_source_source_first;
assign encoder_streamer_sink_sink_last = encoder_source_source_last;
assign encoder_streamer_sink_sink_payload_data = encoder_source_source_payload_data;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_interrupt <= 32'd0;
	hdmi2usbsoc_hdmi2usbsoc_interrupt[1] <= hdmi2usbsoc_hdmi2usbsoc_timer0_irq;
	hdmi2usbsoc_hdmi2usbsoc_interrupt[2] <= hdmi2usbsoc_hdmi2usbsoc_uart_irq;
	hdmi2usbsoc_hdmi2usbsoc_interrupt[4] <= hdmi2usbsoc_hdmi_in0_dma_slot_array_irq;
	hdmi2usbsoc_hdmi2usbsoc_interrupt[5] <= hdmi2usbsoc_hdmi_in1_dma_slot_array_irq;
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_ibus_adr = hdmi2usbsoc_hdmi2usbsoc_i_adr_o[31:2];
assign hdmi2usbsoc_hdmi2usbsoc_dbus_adr = hdmi2usbsoc_hdmi2usbsoc_d_adr_o[31:2];
assign hdmi2usbsoc_hdmi2usbsoc_rom_adr = hdmi2usbsoc_hdmi2usbsoc_rom_bus_adr[12:0];
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_dat_r = hdmi2usbsoc_hdmi2usbsoc_rom_dat_r;

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_sram_we <= 4'd0;
	hdmi2usbsoc_hdmi2usbsoc_sram_we[0] <= (((hdmi2usbsoc_hdmi2usbsoc_sram_bus_cyc & hdmi2usbsoc_hdmi2usbsoc_sram_bus_stb) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_we) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_sel[0]);
	hdmi2usbsoc_hdmi2usbsoc_sram_we[1] <= (((hdmi2usbsoc_hdmi2usbsoc_sram_bus_cyc & hdmi2usbsoc_hdmi2usbsoc_sram_bus_stb) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_we) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_sel[1]);
	hdmi2usbsoc_hdmi2usbsoc_sram_we[2] <= (((hdmi2usbsoc_hdmi2usbsoc_sram_bus_cyc & hdmi2usbsoc_hdmi2usbsoc_sram_bus_stb) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_we) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_sel[2]);
	hdmi2usbsoc_hdmi2usbsoc_sram_we[3] <= (((hdmi2usbsoc_hdmi2usbsoc_sram_bus_cyc & hdmi2usbsoc_hdmi2usbsoc_sram_bus_stb) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_we) & hdmi2usbsoc_hdmi2usbsoc_sram_bus_sel[3]);
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_sram_adr = hdmi2usbsoc_hdmi2usbsoc_sram_bus_adr[11:0];
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_dat_r = hdmi2usbsoc_hdmi2usbsoc_sram_dat_r;
assign hdmi2usbsoc_hdmi2usbsoc_sram_dat_w = hdmi2usbsoc_hdmi2usbsoc_sram_bus_dat_w;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_valid = hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_re;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_payload_data = hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_r;
assign hdmi2usbsoc_hdmi2usbsoc_uart_txfull_status = (~hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_ready);
assign hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_valid = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_valid;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_ready = hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_ready;
assign hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_first = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_first;
assign hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_last = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_last;
assign hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_payload_data = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_trigger = (~hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_ready);
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_valid = hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_valid;
assign hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_ready = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_ready;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_first = hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_first;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_last = hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_last;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_payload_data = hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_payload_data;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rxempty_status = (~hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_valid);
assign hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_w = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_ready = hdmi2usbsoc_hdmi2usbsoc_uart_rx_clear;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_trigger = (~hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_valid);

// synthesis translate_off
reg dummy_d_2;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_uart_tx_clear <= 1'd0;
	if ((hdmi2usbsoc_hdmi2usbsoc_uart_pending_re & hdmi2usbsoc_hdmi2usbsoc_uart_pending_r[0])) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_2 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_3;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_uart_status_w <= 2'd0;
	hdmi2usbsoc_hdmi2usbsoc_uart_status_w[0] <= hdmi2usbsoc_hdmi2usbsoc_uart_tx_status;
	hdmi2usbsoc_hdmi2usbsoc_uart_status_w[1] <= hdmi2usbsoc_hdmi2usbsoc_uart_rx_status;
// synthesis translate_off
	dummy_d_3 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_4;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_uart_rx_clear <= 1'd0;
	if ((hdmi2usbsoc_hdmi2usbsoc_uart_pending_re & hdmi2usbsoc_hdmi2usbsoc_uart_pending_r[1])) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_4 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_5;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_uart_pending_w <= 2'd0;
	hdmi2usbsoc_hdmi2usbsoc_uart_pending_w[0] <= hdmi2usbsoc_hdmi2usbsoc_uart_tx_pending;
	hdmi2usbsoc_hdmi2usbsoc_uart_pending_w[1] <= hdmi2usbsoc_hdmi2usbsoc_uart_rx_pending;
// synthesis translate_off
	dummy_d_5 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_uart_irq = ((hdmi2usbsoc_hdmi2usbsoc_uart_pending_w[0] & hdmi2usbsoc_hdmi2usbsoc_uart_storage[0]) | (hdmi2usbsoc_hdmi2usbsoc_uart_pending_w[1] & hdmi2usbsoc_hdmi2usbsoc_uart_storage[1]));
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_status = hdmi2usbsoc_hdmi2usbsoc_uart_tx_trigger;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_status = hdmi2usbsoc_hdmi2usbsoc_uart_rx_trigger;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_din = {hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_last, hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_first, hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_last, hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_first, hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_ready = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_we = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_valid;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_first = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_first;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_last = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_last;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_valid = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_first = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_last = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_payload_data = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_re = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_source_ready;

// synthesis translate_off
reg dummy_d_6;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_adr <= 4'd0;
	if (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_replace) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_adr <= (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_adr <= hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_6 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_dat_w = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_we = (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_we & (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_writable | hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_replace));
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_do_read = (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_readable & hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_rdport_adr = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_consume;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_dout = hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level != 5'd16);
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_din = {hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_last, hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_first, hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_last, hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_first, hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_ready = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_we = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_valid;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_first = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_first;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_last = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_last;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_valid = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_first = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_last = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_payload_data = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_re = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_source_ready;

// synthesis translate_off
reg dummy_d_7;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_adr <= 4'd0;
	if (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_replace) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_adr <= (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_adr <= hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_7 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_dat_w = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_we = (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_we & (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_writable | hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_replace));
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_do_read = (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_readable & hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_rdport_adr = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_consume;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_dout = hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level != 5'd16);
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi2usbsoc_timer0_zero_trigger = (hdmi2usbsoc_hdmi2usbsoc_timer0_value != 1'd0);
assign hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_status_w = hdmi2usbsoc_hdmi2usbsoc_timer0_zero_status;

// synthesis translate_off
reg dummy_d_8;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi2usbsoc_timer0_zero_clear <= 1'd0;
	if ((hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_re & hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_r)) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_zero_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_8 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_w = hdmi2usbsoc_hdmi2usbsoc_timer0_zero_pending;
assign hdmi2usbsoc_hdmi2usbsoc_timer0_irq = (hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_w & hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage);
assign hdmi2usbsoc_hdmi2usbsoc_timer0_zero_status = hdmi2usbsoc_hdmi2usbsoc_timer0_zero_trigger;
assign por_clk = sys_clk;
assign sdram_full_rd_clk = sdram_full_wr_clk;
assign hdmi2usbsoc_crg_clk4x_rd_strb = hdmi2usbsoc_crg_clk4x_wr_strb;
assign hdmi2usbsoc_git_status = 160'd1286281798330993362540408323602092990343061166500;
assign hdmi2usbsoc_platform_status = 63'd7022356987853668352;
assign hdmi2usbsoc_target_status = 63'd7522257576201122658;
assign hdmi2usbsoc_bus_dat_r = hdmi2usbsoc_sr;

// synthesis translate_off
reg dummy_d_9;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_status <= 1'd0;
	hdmi2usbsoc_o <= 4'd0;
	hdmi2usbsoc_oe <= 1'd0;
	spiflash4x_cs_n <= 1'd0;
	spiflash4x_clk <= 1'd0;
	if (hdmi2usbsoc_bitbang_en_storage) begin
		spiflash4x_clk <= hdmi2usbsoc_bitbang_storage[1];
		spiflash4x_cs_n <= hdmi2usbsoc_bitbang_storage[2];
		if (hdmi2usbsoc_bitbang_storage[3]) begin
			hdmi2usbsoc_oe <= 1'd0;
		end else begin
			hdmi2usbsoc_oe <= 1'd1;
		end
		if (hdmi2usbsoc_bitbang_storage[1]) begin
			hdmi2usbsoc_status <= hdmi2usbsoc_i0[1];
		end
		hdmi2usbsoc_o <= {{3{1'd1}}, hdmi2usbsoc_bitbang_storage[0]};
	end else begin
		spiflash4x_clk <= hdmi2usbsoc_clk;
		spiflash4x_cs_n <= hdmi2usbsoc_cs_n;
		hdmi2usbsoc_o <= hdmi2usbsoc_sr[31:28];
		hdmi2usbsoc_oe <= hdmi2usbsoc_dq_oe;
	end
// synthesis translate_off
	dummy_d_9 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_ddrphy_sdram_half_clk_n = (~sdram_half_clk);
assign hdmi2usbsoc_ddrphy_dqs_t_d0 = (~(hdmi2usbsoc_ddrphy_drive_dqs | hdmi2usbsoc_ddrphy_postamble));
assign hdmi2usbsoc_ddrphy_dqs_t_d1 = (~hdmi2usbsoc_ddrphy_drive_dqs);
assign hdmi2usbsoc_ddrphy_record0_wrdata = hdmi2usbsoc_ddrphy_dfi_p0_wrdata;
assign hdmi2usbsoc_ddrphy_record0_wrdata_mask = hdmi2usbsoc_ddrphy_dfi_p0_wrdata_mask;
assign hdmi2usbsoc_ddrphy_record0_wrdata_en = hdmi2usbsoc_ddrphy_dfi_p0_wrdata_en;
assign hdmi2usbsoc_ddrphy_record0_rddata_en = hdmi2usbsoc_ddrphy_dfi_p0_rddata_en;
assign hdmi2usbsoc_ddrphy_record1_wrdata = hdmi2usbsoc_ddrphy_dfi_p1_wrdata;
assign hdmi2usbsoc_ddrphy_record1_wrdata_mask = hdmi2usbsoc_ddrphy_dfi_p1_wrdata_mask;
assign hdmi2usbsoc_ddrphy_record1_wrdata_en = hdmi2usbsoc_ddrphy_dfi_p1_wrdata_en;
assign hdmi2usbsoc_ddrphy_record1_rddata_en = hdmi2usbsoc_ddrphy_dfi_p1_rddata_en;
assign hdmi2usbsoc_ddrphy_drive_dq_n0 = (~hdmi2usbsoc_ddrphy_drive_dq);
assign hdmi2usbsoc_ddrphy_wrdata_en = (hdmi2usbsoc_ddrphy_record0_wrdata_en | hdmi2usbsoc_ddrphy_record1_wrdata_en);
assign hdmi2usbsoc_ddrphy_drive_dq = hdmi2usbsoc_ddrphy_wrdata_en;
assign hdmi2usbsoc_ddrphy_drive_dqs = hdmi2usbsoc_ddrphy_r_dfi_wrdata_en[1];
assign hdmi2usbsoc_ddrphy_rddata_en = (hdmi2usbsoc_ddrphy_record0_rddata_en | hdmi2usbsoc_ddrphy_record1_rddata_en);
assign hdmi2usbsoc_ddrphy_dfi_p0_rddata = hdmi2usbsoc_ddrphy_record0_rddata;
assign hdmi2usbsoc_ddrphy_dfi_p0_rddata_valid = hdmi2usbsoc_ddrphy_rddata_sr[0];
assign hdmi2usbsoc_ddrphy_dfi_p1_rddata = hdmi2usbsoc_ddrphy_record1_rddata;
assign hdmi2usbsoc_ddrphy_dfi_p1_rddata_valid = hdmi2usbsoc_ddrphy_rddata_sr[0];
assign hdmi2usbsoc_ddrphy_dfi_p0_address = hdmi2usbsoc_sdram_master_p0_address;
assign hdmi2usbsoc_ddrphy_dfi_p0_bank = hdmi2usbsoc_sdram_master_p0_bank;
assign hdmi2usbsoc_ddrphy_dfi_p0_cas_n = hdmi2usbsoc_sdram_master_p0_cas_n;
assign hdmi2usbsoc_ddrphy_dfi_p0_cs_n = hdmi2usbsoc_sdram_master_p0_cs_n;
assign hdmi2usbsoc_ddrphy_dfi_p0_ras_n = hdmi2usbsoc_sdram_master_p0_ras_n;
assign hdmi2usbsoc_ddrphy_dfi_p0_we_n = hdmi2usbsoc_sdram_master_p0_we_n;
assign hdmi2usbsoc_ddrphy_dfi_p0_cke = hdmi2usbsoc_sdram_master_p0_cke;
assign hdmi2usbsoc_ddrphy_dfi_p0_odt = hdmi2usbsoc_sdram_master_p0_odt;
assign hdmi2usbsoc_ddrphy_dfi_p0_reset_n = hdmi2usbsoc_sdram_master_p0_reset_n;
assign hdmi2usbsoc_ddrphy_dfi_p0_wrdata = hdmi2usbsoc_sdram_master_p0_wrdata;
assign hdmi2usbsoc_ddrphy_dfi_p0_wrdata_en = hdmi2usbsoc_sdram_master_p0_wrdata_en;
assign hdmi2usbsoc_ddrphy_dfi_p0_wrdata_mask = hdmi2usbsoc_sdram_master_p0_wrdata_mask;
assign hdmi2usbsoc_ddrphy_dfi_p0_rddata_en = hdmi2usbsoc_sdram_master_p0_rddata_en;
assign hdmi2usbsoc_sdram_master_p0_rddata = hdmi2usbsoc_ddrphy_dfi_p0_rddata;
assign hdmi2usbsoc_sdram_master_p0_rddata_valid = hdmi2usbsoc_ddrphy_dfi_p0_rddata_valid;
assign hdmi2usbsoc_ddrphy_dfi_p1_address = hdmi2usbsoc_sdram_master_p1_address;
assign hdmi2usbsoc_ddrphy_dfi_p1_bank = hdmi2usbsoc_sdram_master_p1_bank;
assign hdmi2usbsoc_ddrphy_dfi_p1_cas_n = hdmi2usbsoc_sdram_master_p1_cas_n;
assign hdmi2usbsoc_ddrphy_dfi_p1_cs_n = hdmi2usbsoc_sdram_master_p1_cs_n;
assign hdmi2usbsoc_ddrphy_dfi_p1_ras_n = hdmi2usbsoc_sdram_master_p1_ras_n;
assign hdmi2usbsoc_ddrphy_dfi_p1_we_n = hdmi2usbsoc_sdram_master_p1_we_n;
assign hdmi2usbsoc_ddrphy_dfi_p1_cke = hdmi2usbsoc_sdram_master_p1_cke;
assign hdmi2usbsoc_ddrphy_dfi_p1_odt = hdmi2usbsoc_sdram_master_p1_odt;
assign hdmi2usbsoc_ddrphy_dfi_p1_reset_n = hdmi2usbsoc_sdram_master_p1_reset_n;
assign hdmi2usbsoc_ddrphy_dfi_p1_wrdata = hdmi2usbsoc_sdram_master_p1_wrdata;
assign hdmi2usbsoc_ddrphy_dfi_p1_wrdata_en = hdmi2usbsoc_sdram_master_p1_wrdata_en;
assign hdmi2usbsoc_ddrphy_dfi_p1_wrdata_mask = hdmi2usbsoc_sdram_master_p1_wrdata_mask;
assign hdmi2usbsoc_ddrphy_dfi_p1_rddata_en = hdmi2usbsoc_sdram_master_p1_rddata_en;
assign hdmi2usbsoc_sdram_master_p1_rddata = hdmi2usbsoc_ddrphy_dfi_p1_rddata;
assign hdmi2usbsoc_sdram_master_p1_rddata_valid = hdmi2usbsoc_ddrphy_dfi_p1_rddata_valid;
assign hdmi2usbsoc_sdram_slave_p0_address = hdmi2usbsoc_sdram_dfi_p0_address;
assign hdmi2usbsoc_sdram_slave_p0_bank = hdmi2usbsoc_sdram_dfi_p0_bank;
assign hdmi2usbsoc_sdram_slave_p0_cas_n = hdmi2usbsoc_sdram_dfi_p0_cas_n;
assign hdmi2usbsoc_sdram_slave_p0_cs_n = hdmi2usbsoc_sdram_dfi_p0_cs_n;
assign hdmi2usbsoc_sdram_slave_p0_ras_n = hdmi2usbsoc_sdram_dfi_p0_ras_n;
assign hdmi2usbsoc_sdram_slave_p0_we_n = hdmi2usbsoc_sdram_dfi_p0_we_n;
assign hdmi2usbsoc_sdram_slave_p0_cke = hdmi2usbsoc_sdram_dfi_p0_cke;
assign hdmi2usbsoc_sdram_slave_p0_odt = hdmi2usbsoc_sdram_dfi_p0_odt;
assign hdmi2usbsoc_sdram_slave_p0_reset_n = hdmi2usbsoc_sdram_dfi_p0_reset_n;
assign hdmi2usbsoc_sdram_slave_p0_wrdata = hdmi2usbsoc_sdram_dfi_p0_wrdata;
assign hdmi2usbsoc_sdram_slave_p0_wrdata_en = hdmi2usbsoc_sdram_dfi_p0_wrdata_en;
assign hdmi2usbsoc_sdram_slave_p0_wrdata_mask = hdmi2usbsoc_sdram_dfi_p0_wrdata_mask;
assign hdmi2usbsoc_sdram_slave_p0_rddata_en = hdmi2usbsoc_sdram_dfi_p0_rddata_en;
assign hdmi2usbsoc_sdram_dfi_p0_rddata = hdmi2usbsoc_sdram_slave_p0_rddata;
assign hdmi2usbsoc_sdram_dfi_p0_rddata_valid = hdmi2usbsoc_sdram_slave_p0_rddata_valid;
assign hdmi2usbsoc_sdram_slave_p1_address = hdmi2usbsoc_sdram_dfi_p1_address;
assign hdmi2usbsoc_sdram_slave_p1_bank = hdmi2usbsoc_sdram_dfi_p1_bank;
assign hdmi2usbsoc_sdram_slave_p1_cas_n = hdmi2usbsoc_sdram_dfi_p1_cas_n;
assign hdmi2usbsoc_sdram_slave_p1_cs_n = hdmi2usbsoc_sdram_dfi_p1_cs_n;
assign hdmi2usbsoc_sdram_slave_p1_ras_n = hdmi2usbsoc_sdram_dfi_p1_ras_n;
assign hdmi2usbsoc_sdram_slave_p1_we_n = hdmi2usbsoc_sdram_dfi_p1_we_n;
assign hdmi2usbsoc_sdram_slave_p1_cke = hdmi2usbsoc_sdram_dfi_p1_cke;
assign hdmi2usbsoc_sdram_slave_p1_odt = hdmi2usbsoc_sdram_dfi_p1_odt;
assign hdmi2usbsoc_sdram_slave_p1_reset_n = hdmi2usbsoc_sdram_dfi_p1_reset_n;
assign hdmi2usbsoc_sdram_slave_p1_wrdata = hdmi2usbsoc_sdram_dfi_p1_wrdata;
assign hdmi2usbsoc_sdram_slave_p1_wrdata_en = hdmi2usbsoc_sdram_dfi_p1_wrdata_en;
assign hdmi2usbsoc_sdram_slave_p1_wrdata_mask = hdmi2usbsoc_sdram_dfi_p1_wrdata_mask;
assign hdmi2usbsoc_sdram_slave_p1_rddata_en = hdmi2usbsoc_sdram_dfi_p1_rddata_en;
assign hdmi2usbsoc_sdram_dfi_p1_rddata = hdmi2usbsoc_sdram_slave_p1_rddata;
assign hdmi2usbsoc_sdram_dfi_p1_rddata_valid = hdmi2usbsoc_sdram_slave_p1_rddata_valid;

// synthesis translate_off
reg dummy_d_10;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_inti_p0_rddata <= 32'd0;
	hdmi2usbsoc_sdram_inti_p0_rddata_valid <= 1'd0;
	hdmi2usbsoc_sdram_inti_p1_rddata <= 32'd0;
	hdmi2usbsoc_sdram_inti_p1_rddata_valid <= 1'd0;
	hdmi2usbsoc_sdram_slave_p0_rddata <= 32'd0;
	hdmi2usbsoc_sdram_slave_p0_rddata_valid <= 1'd0;
	hdmi2usbsoc_sdram_slave_p1_rddata <= 32'd0;
	hdmi2usbsoc_sdram_slave_p1_rddata_valid <= 1'd0;
	hdmi2usbsoc_sdram_master_p0_address <= 13'd0;
	hdmi2usbsoc_sdram_master_p0_bank <= 3'd0;
	hdmi2usbsoc_sdram_master_p0_cas_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p0_cs_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p0_ras_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p0_we_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p0_cke <= 1'd0;
	hdmi2usbsoc_sdram_master_p0_odt <= 1'd0;
	hdmi2usbsoc_sdram_master_p0_reset_n <= 1'd0;
	hdmi2usbsoc_sdram_master_p0_wrdata <= 32'd0;
	hdmi2usbsoc_sdram_master_p0_wrdata_en <= 1'd0;
	hdmi2usbsoc_sdram_master_p0_wrdata_mask <= 4'd0;
	hdmi2usbsoc_sdram_master_p0_rddata_en <= 1'd0;
	hdmi2usbsoc_sdram_master_p1_address <= 13'd0;
	hdmi2usbsoc_sdram_master_p1_bank <= 3'd0;
	hdmi2usbsoc_sdram_master_p1_cas_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p1_cs_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p1_ras_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p1_we_n <= 1'd1;
	hdmi2usbsoc_sdram_master_p1_cke <= 1'd0;
	hdmi2usbsoc_sdram_master_p1_odt <= 1'd0;
	hdmi2usbsoc_sdram_master_p1_reset_n <= 1'd0;
	hdmi2usbsoc_sdram_master_p1_wrdata <= 32'd0;
	hdmi2usbsoc_sdram_master_p1_wrdata_en <= 1'd0;
	hdmi2usbsoc_sdram_master_p1_wrdata_mask <= 4'd0;
	hdmi2usbsoc_sdram_master_p1_rddata_en <= 1'd0;
	if (hdmi2usbsoc_sdram_storage[0]) begin
		hdmi2usbsoc_sdram_master_p0_address <= hdmi2usbsoc_sdram_slave_p0_address;
		hdmi2usbsoc_sdram_master_p0_bank <= hdmi2usbsoc_sdram_slave_p0_bank;
		hdmi2usbsoc_sdram_master_p0_cas_n <= hdmi2usbsoc_sdram_slave_p0_cas_n;
		hdmi2usbsoc_sdram_master_p0_cs_n <= hdmi2usbsoc_sdram_slave_p0_cs_n;
		hdmi2usbsoc_sdram_master_p0_ras_n <= hdmi2usbsoc_sdram_slave_p0_ras_n;
		hdmi2usbsoc_sdram_master_p0_we_n <= hdmi2usbsoc_sdram_slave_p0_we_n;
		hdmi2usbsoc_sdram_master_p0_cke <= hdmi2usbsoc_sdram_slave_p0_cke;
		hdmi2usbsoc_sdram_master_p0_odt <= hdmi2usbsoc_sdram_slave_p0_odt;
		hdmi2usbsoc_sdram_master_p0_reset_n <= hdmi2usbsoc_sdram_slave_p0_reset_n;
		hdmi2usbsoc_sdram_master_p0_wrdata <= hdmi2usbsoc_sdram_slave_p0_wrdata;
		hdmi2usbsoc_sdram_master_p0_wrdata_en <= hdmi2usbsoc_sdram_slave_p0_wrdata_en;
		hdmi2usbsoc_sdram_master_p0_wrdata_mask <= hdmi2usbsoc_sdram_slave_p0_wrdata_mask;
		hdmi2usbsoc_sdram_master_p0_rddata_en <= hdmi2usbsoc_sdram_slave_p0_rddata_en;
		hdmi2usbsoc_sdram_slave_p0_rddata <= hdmi2usbsoc_sdram_master_p0_rddata;
		hdmi2usbsoc_sdram_slave_p0_rddata_valid <= hdmi2usbsoc_sdram_master_p0_rddata_valid;
		hdmi2usbsoc_sdram_master_p1_address <= hdmi2usbsoc_sdram_slave_p1_address;
		hdmi2usbsoc_sdram_master_p1_bank <= hdmi2usbsoc_sdram_slave_p1_bank;
		hdmi2usbsoc_sdram_master_p1_cas_n <= hdmi2usbsoc_sdram_slave_p1_cas_n;
		hdmi2usbsoc_sdram_master_p1_cs_n <= hdmi2usbsoc_sdram_slave_p1_cs_n;
		hdmi2usbsoc_sdram_master_p1_ras_n <= hdmi2usbsoc_sdram_slave_p1_ras_n;
		hdmi2usbsoc_sdram_master_p1_we_n <= hdmi2usbsoc_sdram_slave_p1_we_n;
		hdmi2usbsoc_sdram_master_p1_cke <= hdmi2usbsoc_sdram_slave_p1_cke;
		hdmi2usbsoc_sdram_master_p1_odt <= hdmi2usbsoc_sdram_slave_p1_odt;
		hdmi2usbsoc_sdram_master_p1_reset_n <= hdmi2usbsoc_sdram_slave_p1_reset_n;
		hdmi2usbsoc_sdram_master_p1_wrdata <= hdmi2usbsoc_sdram_slave_p1_wrdata;
		hdmi2usbsoc_sdram_master_p1_wrdata_en <= hdmi2usbsoc_sdram_slave_p1_wrdata_en;
		hdmi2usbsoc_sdram_master_p1_wrdata_mask <= hdmi2usbsoc_sdram_slave_p1_wrdata_mask;
		hdmi2usbsoc_sdram_master_p1_rddata_en <= hdmi2usbsoc_sdram_slave_p1_rddata_en;
		hdmi2usbsoc_sdram_slave_p1_rddata <= hdmi2usbsoc_sdram_master_p1_rddata;
		hdmi2usbsoc_sdram_slave_p1_rddata_valid <= hdmi2usbsoc_sdram_master_p1_rddata_valid;
	end else begin
		hdmi2usbsoc_sdram_master_p0_address <= hdmi2usbsoc_sdram_inti_p0_address;
		hdmi2usbsoc_sdram_master_p0_bank <= hdmi2usbsoc_sdram_inti_p0_bank;
		hdmi2usbsoc_sdram_master_p0_cas_n <= hdmi2usbsoc_sdram_inti_p0_cas_n;
		hdmi2usbsoc_sdram_master_p0_cs_n <= hdmi2usbsoc_sdram_inti_p0_cs_n;
		hdmi2usbsoc_sdram_master_p0_ras_n <= hdmi2usbsoc_sdram_inti_p0_ras_n;
		hdmi2usbsoc_sdram_master_p0_we_n <= hdmi2usbsoc_sdram_inti_p0_we_n;
		hdmi2usbsoc_sdram_master_p0_cke <= hdmi2usbsoc_sdram_inti_p0_cke;
		hdmi2usbsoc_sdram_master_p0_odt <= hdmi2usbsoc_sdram_inti_p0_odt;
		hdmi2usbsoc_sdram_master_p0_reset_n <= hdmi2usbsoc_sdram_inti_p0_reset_n;
		hdmi2usbsoc_sdram_master_p0_wrdata <= hdmi2usbsoc_sdram_inti_p0_wrdata;
		hdmi2usbsoc_sdram_master_p0_wrdata_en <= hdmi2usbsoc_sdram_inti_p0_wrdata_en;
		hdmi2usbsoc_sdram_master_p0_wrdata_mask <= hdmi2usbsoc_sdram_inti_p0_wrdata_mask;
		hdmi2usbsoc_sdram_master_p0_rddata_en <= hdmi2usbsoc_sdram_inti_p0_rddata_en;
		hdmi2usbsoc_sdram_inti_p0_rddata <= hdmi2usbsoc_sdram_master_p0_rddata;
		hdmi2usbsoc_sdram_inti_p0_rddata_valid <= hdmi2usbsoc_sdram_master_p0_rddata_valid;
		hdmi2usbsoc_sdram_master_p1_address <= hdmi2usbsoc_sdram_inti_p1_address;
		hdmi2usbsoc_sdram_master_p1_bank <= hdmi2usbsoc_sdram_inti_p1_bank;
		hdmi2usbsoc_sdram_master_p1_cas_n <= hdmi2usbsoc_sdram_inti_p1_cas_n;
		hdmi2usbsoc_sdram_master_p1_cs_n <= hdmi2usbsoc_sdram_inti_p1_cs_n;
		hdmi2usbsoc_sdram_master_p1_ras_n <= hdmi2usbsoc_sdram_inti_p1_ras_n;
		hdmi2usbsoc_sdram_master_p1_we_n <= hdmi2usbsoc_sdram_inti_p1_we_n;
		hdmi2usbsoc_sdram_master_p1_cke <= hdmi2usbsoc_sdram_inti_p1_cke;
		hdmi2usbsoc_sdram_master_p1_odt <= hdmi2usbsoc_sdram_inti_p1_odt;
		hdmi2usbsoc_sdram_master_p1_reset_n <= hdmi2usbsoc_sdram_inti_p1_reset_n;
		hdmi2usbsoc_sdram_master_p1_wrdata <= hdmi2usbsoc_sdram_inti_p1_wrdata;
		hdmi2usbsoc_sdram_master_p1_wrdata_en <= hdmi2usbsoc_sdram_inti_p1_wrdata_en;
		hdmi2usbsoc_sdram_master_p1_wrdata_mask <= hdmi2usbsoc_sdram_inti_p1_wrdata_mask;
		hdmi2usbsoc_sdram_master_p1_rddata_en <= hdmi2usbsoc_sdram_inti_p1_rddata_en;
		hdmi2usbsoc_sdram_inti_p1_rddata <= hdmi2usbsoc_sdram_master_p1_rddata;
		hdmi2usbsoc_sdram_inti_p1_rddata_valid <= hdmi2usbsoc_sdram_master_p1_rddata_valid;
	end
// synthesis translate_off
	dummy_d_10 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_inti_p0_cke = hdmi2usbsoc_sdram_storage[1];
assign hdmi2usbsoc_sdram_inti_p1_cke = hdmi2usbsoc_sdram_storage[1];
assign hdmi2usbsoc_sdram_inti_p0_odt = hdmi2usbsoc_sdram_storage[2];
assign hdmi2usbsoc_sdram_inti_p1_odt = hdmi2usbsoc_sdram_storage[2];
assign hdmi2usbsoc_sdram_inti_p0_reset_n = hdmi2usbsoc_sdram_storage[3];
assign hdmi2usbsoc_sdram_inti_p1_reset_n = hdmi2usbsoc_sdram_storage[3];

// synthesis translate_off
reg dummy_d_11;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_inti_p0_cas_n <= 1'd1;
	hdmi2usbsoc_sdram_inti_p0_cs_n <= 1'd1;
	hdmi2usbsoc_sdram_inti_p0_ras_n <= 1'd1;
	hdmi2usbsoc_sdram_inti_p0_we_n <= 1'd1;
	if (hdmi2usbsoc_sdram_phaseinjector0_command_issue_re) begin
		hdmi2usbsoc_sdram_inti_p0_cs_n <= (~hdmi2usbsoc_sdram_phaseinjector0_command_storage[0]);
		hdmi2usbsoc_sdram_inti_p0_we_n <= (~hdmi2usbsoc_sdram_phaseinjector0_command_storage[1]);
		hdmi2usbsoc_sdram_inti_p0_cas_n <= (~hdmi2usbsoc_sdram_phaseinjector0_command_storage[2]);
		hdmi2usbsoc_sdram_inti_p0_ras_n <= (~hdmi2usbsoc_sdram_phaseinjector0_command_storage[3]);
	end else begin
		hdmi2usbsoc_sdram_inti_p0_cs_n <= 1'd1;
		hdmi2usbsoc_sdram_inti_p0_we_n <= 1'd1;
		hdmi2usbsoc_sdram_inti_p0_cas_n <= 1'd1;
		hdmi2usbsoc_sdram_inti_p0_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_11 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_inti_p0_address = hdmi2usbsoc_sdram_phaseinjector0_address_storage;
assign hdmi2usbsoc_sdram_inti_p0_bank = hdmi2usbsoc_sdram_phaseinjector0_baddress_storage;
assign hdmi2usbsoc_sdram_inti_p0_wrdata_en = (hdmi2usbsoc_sdram_phaseinjector0_command_issue_re & hdmi2usbsoc_sdram_phaseinjector0_command_storage[4]);
assign hdmi2usbsoc_sdram_inti_p0_rddata_en = (hdmi2usbsoc_sdram_phaseinjector0_command_issue_re & hdmi2usbsoc_sdram_phaseinjector0_command_storage[5]);
assign hdmi2usbsoc_sdram_inti_p0_wrdata = hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage;
assign hdmi2usbsoc_sdram_inti_p0_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_12;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_inti_p1_cs_n <= 1'd1;
	hdmi2usbsoc_sdram_inti_p1_ras_n <= 1'd1;
	hdmi2usbsoc_sdram_inti_p1_we_n <= 1'd1;
	hdmi2usbsoc_sdram_inti_p1_cas_n <= 1'd1;
	if (hdmi2usbsoc_sdram_phaseinjector1_command_issue_re) begin
		hdmi2usbsoc_sdram_inti_p1_cs_n <= (~hdmi2usbsoc_sdram_phaseinjector1_command_storage[0]);
		hdmi2usbsoc_sdram_inti_p1_we_n <= (~hdmi2usbsoc_sdram_phaseinjector1_command_storage[1]);
		hdmi2usbsoc_sdram_inti_p1_cas_n <= (~hdmi2usbsoc_sdram_phaseinjector1_command_storage[2]);
		hdmi2usbsoc_sdram_inti_p1_ras_n <= (~hdmi2usbsoc_sdram_phaseinjector1_command_storage[3]);
	end else begin
		hdmi2usbsoc_sdram_inti_p1_cs_n <= 1'd1;
		hdmi2usbsoc_sdram_inti_p1_we_n <= 1'd1;
		hdmi2usbsoc_sdram_inti_p1_cas_n <= 1'd1;
		hdmi2usbsoc_sdram_inti_p1_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_12 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_inti_p1_address = hdmi2usbsoc_sdram_phaseinjector1_address_storage;
assign hdmi2usbsoc_sdram_inti_p1_bank = hdmi2usbsoc_sdram_phaseinjector1_baddress_storage;
assign hdmi2usbsoc_sdram_inti_p1_wrdata_en = (hdmi2usbsoc_sdram_phaseinjector1_command_issue_re & hdmi2usbsoc_sdram_phaseinjector1_command_storage[4]);
assign hdmi2usbsoc_sdram_inti_p1_rddata_en = (hdmi2usbsoc_sdram_phaseinjector1_command_issue_re & hdmi2usbsoc_sdram_phaseinjector1_command_storage[5]);
assign hdmi2usbsoc_sdram_inti_p1_wrdata = hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage;
assign hdmi2usbsoc_sdram_inti_p1_wrdata_mask = 1'd0;
assign hdmi2usbsoc_sdram_bankmachine0_req_valid = hdmi2usbsoc_sdram_interface_bank0_valid;
assign hdmi2usbsoc_sdram_interface_bank0_ready = hdmi2usbsoc_sdram_bankmachine0_req_ready;
assign hdmi2usbsoc_sdram_bankmachine0_req_we = hdmi2usbsoc_sdram_interface_bank0_we;
assign hdmi2usbsoc_sdram_bankmachine0_req_adr = hdmi2usbsoc_sdram_interface_bank0_adr;
assign hdmi2usbsoc_sdram_interface_bank0_lock = hdmi2usbsoc_sdram_bankmachine0_req_lock;
assign hdmi2usbsoc_sdram_interface_bank0_wdata_ready = hdmi2usbsoc_sdram_bankmachine0_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank0_rdata_valid = hdmi2usbsoc_sdram_bankmachine0_req_rdata_valid;
assign hdmi2usbsoc_sdram_bankmachine1_req_valid = hdmi2usbsoc_sdram_interface_bank1_valid;
assign hdmi2usbsoc_sdram_interface_bank1_ready = hdmi2usbsoc_sdram_bankmachine1_req_ready;
assign hdmi2usbsoc_sdram_bankmachine1_req_we = hdmi2usbsoc_sdram_interface_bank1_we;
assign hdmi2usbsoc_sdram_bankmachine1_req_adr = hdmi2usbsoc_sdram_interface_bank1_adr;
assign hdmi2usbsoc_sdram_interface_bank1_lock = hdmi2usbsoc_sdram_bankmachine1_req_lock;
assign hdmi2usbsoc_sdram_interface_bank1_wdata_ready = hdmi2usbsoc_sdram_bankmachine1_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank1_rdata_valid = hdmi2usbsoc_sdram_bankmachine1_req_rdata_valid;
assign hdmi2usbsoc_sdram_bankmachine2_req_valid = hdmi2usbsoc_sdram_interface_bank2_valid;
assign hdmi2usbsoc_sdram_interface_bank2_ready = hdmi2usbsoc_sdram_bankmachine2_req_ready;
assign hdmi2usbsoc_sdram_bankmachine2_req_we = hdmi2usbsoc_sdram_interface_bank2_we;
assign hdmi2usbsoc_sdram_bankmachine2_req_adr = hdmi2usbsoc_sdram_interface_bank2_adr;
assign hdmi2usbsoc_sdram_interface_bank2_lock = hdmi2usbsoc_sdram_bankmachine2_req_lock;
assign hdmi2usbsoc_sdram_interface_bank2_wdata_ready = hdmi2usbsoc_sdram_bankmachine2_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank2_rdata_valid = hdmi2usbsoc_sdram_bankmachine2_req_rdata_valid;
assign hdmi2usbsoc_sdram_bankmachine3_req_valid = hdmi2usbsoc_sdram_interface_bank3_valid;
assign hdmi2usbsoc_sdram_interface_bank3_ready = hdmi2usbsoc_sdram_bankmachine3_req_ready;
assign hdmi2usbsoc_sdram_bankmachine3_req_we = hdmi2usbsoc_sdram_interface_bank3_we;
assign hdmi2usbsoc_sdram_bankmachine3_req_adr = hdmi2usbsoc_sdram_interface_bank3_adr;
assign hdmi2usbsoc_sdram_interface_bank3_lock = hdmi2usbsoc_sdram_bankmachine3_req_lock;
assign hdmi2usbsoc_sdram_interface_bank3_wdata_ready = hdmi2usbsoc_sdram_bankmachine3_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank3_rdata_valid = hdmi2usbsoc_sdram_bankmachine3_req_rdata_valid;
assign hdmi2usbsoc_sdram_bankmachine4_req_valid = hdmi2usbsoc_sdram_interface_bank4_valid;
assign hdmi2usbsoc_sdram_interface_bank4_ready = hdmi2usbsoc_sdram_bankmachine4_req_ready;
assign hdmi2usbsoc_sdram_bankmachine4_req_we = hdmi2usbsoc_sdram_interface_bank4_we;
assign hdmi2usbsoc_sdram_bankmachine4_req_adr = hdmi2usbsoc_sdram_interface_bank4_adr;
assign hdmi2usbsoc_sdram_interface_bank4_lock = hdmi2usbsoc_sdram_bankmachine4_req_lock;
assign hdmi2usbsoc_sdram_interface_bank4_wdata_ready = hdmi2usbsoc_sdram_bankmachine4_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank4_rdata_valid = hdmi2usbsoc_sdram_bankmachine4_req_rdata_valid;
assign hdmi2usbsoc_sdram_bankmachine5_req_valid = hdmi2usbsoc_sdram_interface_bank5_valid;
assign hdmi2usbsoc_sdram_interface_bank5_ready = hdmi2usbsoc_sdram_bankmachine5_req_ready;
assign hdmi2usbsoc_sdram_bankmachine5_req_we = hdmi2usbsoc_sdram_interface_bank5_we;
assign hdmi2usbsoc_sdram_bankmachine5_req_adr = hdmi2usbsoc_sdram_interface_bank5_adr;
assign hdmi2usbsoc_sdram_interface_bank5_lock = hdmi2usbsoc_sdram_bankmachine5_req_lock;
assign hdmi2usbsoc_sdram_interface_bank5_wdata_ready = hdmi2usbsoc_sdram_bankmachine5_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank5_rdata_valid = hdmi2usbsoc_sdram_bankmachine5_req_rdata_valid;
assign hdmi2usbsoc_sdram_bankmachine6_req_valid = hdmi2usbsoc_sdram_interface_bank6_valid;
assign hdmi2usbsoc_sdram_interface_bank6_ready = hdmi2usbsoc_sdram_bankmachine6_req_ready;
assign hdmi2usbsoc_sdram_bankmachine6_req_we = hdmi2usbsoc_sdram_interface_bank6_we;
assign hdmi2usbsoc_sdram_bankmachine6_req_adr = hdmi2usbsoc_sdram_interface_bank6_adr;
assign hdmi2usbsoc_sdram_interface_bank6_lock = hdmi2usbsoc_sdram_bankmachine6_req_lock;
assign hdmi2usbsoc_sdram_interface_bank6_wdata_ready = hdmi2usbsoc_sdram_bankmachine6_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank6_rdata_valid = hdmi2usbsoc_sdram_bankmachine6_req_rdata_valid;
assign hdmi2usbsoc_sdram_bankmachine7_req_valid = hdmi2usbsoc_sdram_interface_bank7_valid;
assign hdmi2usbsoc_sdram_interface_bank7_ready = hdmi2usbsoc_sdram_bankmachine7_req_ready;
assign hdmi2usbsoc_sdram_bankmachine7_req_we = hdmi2usbsoc_sdram_interface_bank7_we;
assign hdmi2usbsoc_sdram_bankmachine7_req_adr = hdmi2usbsoc_sdram_interface_bank7_adr;
assign hdmi2usbsoc_sdram_interface_bank7_lock = hdmi2usbsoc_sdram_bankmachine7_req_lock;
assign hdmi2usbsoc_sdram_interface_bank7_wdata_ready = hdmi2usbsoc_sdram_bankmachine7_req_wdata_ready;
assign hdmi2usbsoc_sdram_interface_bank7_rdata_valid = hdmi2usbsoc_sdram_bankmachine7_req_rdata_valid;
assign hdmi2usbsoc_sdram_wait = (1'd1 & (~hdmi2usbsoc_sdram_done));
assign hdmi2usbsoc_sdram_done = (hdmi2usbsoc_sdram_count == 1'd0);

// synthesis translate_off
reg dummy_d_13;
// synthesis translate_on
always @(*) begin
	controllerinjector_refresher_next_state <= 2'd0;
	hdmi2usbsoc_sdram_cmd_valid <= 1'd0;
	hdmi2usbsoc_sdram_cmd_last <= 1'd0;
	hdmi2usbsoc_sdram_seq_start <= 1'd0;
	controllerinjector_refresher_next_state <= controllerinjector_refresher_state;
	case (controllerinjector_refresher_state)
		1'd1: begin
			hdmi2usbsoc_sdram_cmd_valid <= 1'd1;
			if (hdmi2usbsoc_sdram_cmd_ready) begin
				hdmi2usbsoc_sdram_seq_start <= 1'd1;
				controllerinjector_refresher_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (hdmi2usbsoc_sdram_seq_done) begin
				hdmi2usbsoc_sdram_cmd_last <= 1'd1;
				controllerinjector_refresher_next_state <= 1'd0;
			end else begin
				hdmi2usbsoc_sdram_cmd_valid <= 1'd1;
			end
		end
		default: begin
			if (hdmi2usbsoc_sdram_done) begin
				controllerinjector_refresher_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_13 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine0_sink_valid = hdmi2usbsoc_sdram_bankmachine0_req_valid;
assign hdmi2usbsoc_sdram_bankmachine0_req_ready = hdmi2usbsoc_sdram_bankmachine0_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine0_sink_payload_we = hdmi2usbsoc_sdram_bankmachine0_req_we;
assign hdmi2usbsoc_sdram_bankmachine0_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine0_req_adr;
assign hdmi2usbsoc_sdram_bankmachine0_source_ready = (hdmi2usbsoc_sdram_bankmachine0_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine0_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine0_req_lock = hdmi2usbsoc_sdram_bankmachine0_source_valid;
assign hdmi2usbsoc_sdram_bankmachine0_hit = (hdmi2usbsoc_sdram_bankmachine0_openrow == hdmi2usbsoc_sdram_bankmachine0_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ba = 1'd0;

// synthesis translate_off
reg dummy_d_14;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine0_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine0_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine0_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine0_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine0_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine0_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_14 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine0_wait = (~((hdmi2usbsoc_sdram_bankmachine0_cmd_valid & hdmi2usbsoc_sdram_bankmachine0_cmd_ready) & hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine0_syncfifo0_din = {hdmi2usbsoc_sdram_bankmachine0_fifo_in_last, hdmi2usbsoc_sdram_bankmachine0_fifo_in_first, hdmi2usbsoc_sdram_bankmachine0_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine0_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine0_fifo_out_last, hdmi2usbsoc_sdram_bankmachine0_fifo_out_first, hdmi2usbsoc_sdram_bankmachine0_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine0_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine0_syncfifo0_dout;
assign hdmi2usbsoc_sdram_bankmachine0_sink_ready = hdmi2usbsoc_sdram_bankmachine0_syncfifo0_writable;
assign hdmi2usbsoc_sdram_bankmachine0_syncfifo0_we = hdmi2usbsoc_sdram_bankmachine0_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine0_fifo_in_first = hdmi2usbsoc_sdram_bankmachine0_sink_first;
assign hdmi2usbsoc_sdram_bankmachine0_fifo_in_last = hdmi2usbsoc_sdram_bankmachine0_sink_last;
assign hdmi2usbsoc_sdram_bankmachine0_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine0_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine0_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine0_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine0_source_valid = hdmi2usbsoc_sdram_bankmachine0_syncfifo0_readable;
assign hdmi2usbsoc_sdram_bankmachine0_source_first = hdmi2usbsoc_sdram_bankmachine0_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine0_source_last = hdmi2usbsoc_sdram_bankmachine0_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine0_source_payload_we = hdmi2usbsoc_sdram_bankmachine0_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine0_source_payload_adr = hdmi2usbsoc_sdram_bankmachine0_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine0_syncfifo0_re = hdmi2usbsoc_sdram_bankmachine0_source_ready;

// synthesis translate_off
reg dummy_d_15;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine0_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine0_replace) begin
		hdmi2usbsoc_sdram_bankmachine0_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine0_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine0_wrport_adr <= hdmi2usbsoc_sdram_bankmachine0_produce;
	end
// synthesis translate_off
	dummy_d_15 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine0_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine0_syncfifo0_din;
assign hdmi2usbsoc_sdram_bankmachine0_wrport_we = (hdmi2usbsoc_sdram_bankmachine0_syncfifo0_we & (hdmi2usbsoc_sdram_bankmachine0_syncfifo0_writable | hdmi2usbsoc_sdram_bankmachine0_replace));
assign hdmi2usbsoc_sdram_bankmachine0_do_read = (hdmi2usbsoc_sdram_bankmachine0_syncfifo0_readable & hdmi2usbsoc_sdram_bankmachine0_syncfifo0_re);
assign hdmi2usbsoc_sdram_bankmachine0_rdport_adr = hdmi2usbsoc_sdram_bankmachine0_consume;
assign hdmi2usbsoc_sdram_bankmachine0_syncfifo0_dout = hdmi2usbsoc_sdram_bankmachine0_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine0_syncfifo0_writable = (hdmi2usbsoc_sdram_bankmachine0_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine0_syncfifo0_readable = (hdmi2usbsoc_sdram_bankmachine0_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine0_done = (hdmi2usbsoc_sdram_bankmachine0_count == 1'd0);

// synthesis translate_off
reg dummy_d_16;
// synthesis translate_on
always @(*) begin
	controllerinjector_bankmachine0_next_state <= 3'd0;
	hdmi2usbsoc_sdram_bankmachine0_req_wdata_ready <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_req_rdata_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_cmd_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_sel_row_adr <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd0;
	controllerinjector_bankmachine0_next_state <= controllerinjector_bankmachine0_state;
	case (controllerinjector_bankmachine0_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine0_done) begin
				hdmi2usbsoc_sdram_bankmachine0_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine0_cmd_ready) begin
					controllerinjector_bankmachine0_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine0_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine0_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine0_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine0_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine0_cmd_ready) begin
				controllerinjector_bankmachine0_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine0_done) begin
				hdmi2usbsoc_sdram_bankmachine0_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine0_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine0_refresh_req)) begin
				controllerinjector_bankmachine0_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine0_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine0_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine0_refresh_req) begin
				controllerinjector_bankmachine0_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine0_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine0_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine0_hit) begin
							hdmi2usbsoc_sdram_bankmachine0_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine0_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine0_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine0_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine0_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine0_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine0_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine0_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine0_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_16 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine1_sink_valid = hdmi2usbsoc_sdram_bankmachine1_req_valid;
assign hdmi2usbsoc_sdram_bankmachine1_req_ready = hdmi2usbsoc_sdram_bankmachine1_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine1_sink_payload_we = hdmi2usbsoc_sdram_bankmachine1_req_we;
assign hdmi2usbsoc_sdram_bankmachine1_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine1_req_adr;
assign hdmi2usbsoc_sdram_bankmachine1_source_ready = (hdmi2usbsoc_sdram_bankmachine1_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine1_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine1_req_lock = hdmi2usbsoc_sdram_bankmachine1_source_valid;
assign hdmi2usbsoc_sdram_bankmachine1_hit = (hdmi2usbsoc_sdram_bankmachine1_openrow == hdmi2usbsoc_sdram_bankmachine1_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ba = 1'd1;

// synthesis translate_off
reg dummy_d_17;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine1_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine1_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine1_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine1_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine1_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine1_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_17 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine1_wait = (~((hdmi2usbsoc_sdram_bankmachine1_cmd_valid & hdmi2usbsoc_sdram_bankmachine1_cmd_ready) & hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine1_syncfifo1_din = {hdmi2usbsoc_sdram_bankmachine1_fifo_in_last, hdmi2usbsoc_sdram_bankmachine1_fifo_in_first, hdmi2usbsoc_sdram_bankmachine1_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine1_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine1_fifo_out_last, hdmi2usbsoc_sdram_bankmachine1_fifo_out_first, hdmi2usbsoc_sdram_bankmachine1_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine1_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine1_syncfifo1_dout;
assign hdmi2usbsoc_sdram_bankmachine1_sink_ready = hdmi2usbsoc_sdram_bankmachine1_syncfifo1_writable;
assign hdmi2usbsoc_sdram_bankmachine1_syncfifo1_we = hdmi2usbsoc_sdram_bankmachine1_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine1_fifo_in_first = hdmi2usbsoc_sdram_bankmachine1_sink_first;
assign hdmi2usbsoc_sdram_bankmachine1_fifo_in_last = hdmi2usbsoc_sdram_bankmachine1_sink_last;
assign hdmi2usbsoc_sdram_bankmachine1_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine1_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine1_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine1_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine1_source_valid = hdmi2usbsoc_sdram_bankmachine1_syncfifo1_readable;
assign hdmi2usbsoc_sdram_bankmachine1_source_first = hdmi2usbsoc_sdram_bankmachine1_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine1_source_last = hdmi2usbsoc_sdram_bankmachine1_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine1_source_payload_we = hdmi2usbsoc_sdram_bankmachine1_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine1_source_payload_adr = hdmi2usbsoc_sdram_bankmachine1_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine1_syncfifo1_re = hdmi2usbsoc_sdram_bankmachine1_source_ready;

// synthesis translate_off
reg dummy_d_18;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine1_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine1_replace) begin
		hdmi2usbsoc_sdram_bankmachine1_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine1_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine1_wrport_adr <= hdmi2usbsoc_sdram_bankmachine1_produce;
	end
// synthesis translate_off
	dummy_d_18 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine1_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine1_syncfifo1_din;
assign hdmi2usbsoc_sdram_bankmachine1_wrport_we = (hdmi2usbsoc_sdram_bankmachine1_syncfifo1_we & (hdmi2usbsoc_sdram_bankmachine1_syncfifo1_writable | hdmi2usbsoc_sdram_bankmachine1_replace));
assign hdmi2usbsoc_sdram_bankmachine1_do_read = (hdmi2usbsoc_sdram_bankmachine1_syncfifo1_readable & hdmi2usbsoc_sdram_bankmachine1_syncfifo1_re);
assign hdmi2usbsoc_sdram_bankmachine1_rdport_adr = hdmi2usbsoc_sdram_bankmachine1_consume;
assign hdmi2usbsoc_sdram_bankmachine1_syncfifo1_dout = hdmi2usbsoc_sdram_bankmachine1_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine1_syncfifo1_writable = (hdmi2usbsoc_sdram_bankmachine1_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine1_syncfifo1_readable = (hdmi2usbsoc_sdram_bankmachine1_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine1_done = (hdmi2usbsoc_sdram_bankmachine1_count == 1'd0);

// synthesis translate_off
reg dummy_d_19;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_req_wdata_ready <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_req_rdata_valid <= 1'd0;
	controllerinjector_bankmachine1_next_state <= 3'd0;
	hdmi2usbsoc_sdram_bankmachine1_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_cmd_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine1_sel_row_adr <= 1'd0;
	controllerinjector_bankmachine1_next_state <= controllerinjector_bankmachine1_state;
	case (controllerinjector_bankmachine1_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine1_done) begin
				hdmi2usbsoc_sdram_bankmachine1_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine1_cmd_ready) begin
					controllerinjector_bankmachine1_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine1_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine1_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine1_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine1_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine1_cmd_ready) begin
				controllerinjector_bankmachine1_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine1_done) begin
				hdmi2usbsoc_sdram_bankmachine1_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine1_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine1_refresh_req)) begin
				controllerinjector_bankmachine1_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine1_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine1_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine1_refresh_req) begin
				controllerinjector_bankmachine1_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine1_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine1_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine1_hit) begin
							hdmi2usbsoc_sdram_bankmachine1_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine1_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine1_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine1_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine1_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine1_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine1_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine1_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine1_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_19 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine2_sink_valid = hdmi2usbsoc_sdram_bankmachine2_req_valid;
assign hdmi2usbsoc_sdram_bankmachine2_req_ready = hdmi2usbsoc_sdram_bankmachine2_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine2_sink_payload_we = hdmi2usbsoc_sdram_bankmachine2_req_we;
assign hdmi2usbsoc_sdram_bankmachine2_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine2_req_adr;
assign hdmi2usbsoc_sdram_bankmachine2_source_ready = (hdmi2usbsoc_sdram_bankmachine2_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine2_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine2_req_lock = hdmi2usbsoc_sdram_bankmachine2_source_valid;
assign hdmi2usbsoc_sdram_bankmachine2_hit = (hdmi2usbsoc_sdram_bankmachine2_openrow == hdmi2usbsoc_sdram_bankmachine2_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ba = 2'd2;

// synthesis translate_off
reg dummy_d_20;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine2_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine2_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine2_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine2_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine2_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine2_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_20 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine2_wait = (~((hdmi2usbsoc_sdram_bankmachine2_cmd_valid & hdmi2usbsoc_sdram_bankmachine2_cmd_ready) & hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine2_syncfifo2_din = {hdmi2usbsoc_sdram_bankmachine2_fifo_in_last, hdmi2usbsoc_sdram_bankmachine2_fifo_in_first, hdmi2usbsoc_sdram_bankmachine2_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine2_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine2_fifo_out_last, hdmi2usbsoc_sdram_bankmachine2_fifo_out_first, hdmi2usbsoc_sdram_bankmachine2_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine2_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine2_syncfifo2_dout;
assign hdmi2usbsoc_sdram_bankmachine2_sink_ready = hdmi2usbsoc_sdram_bankmachine2_syncfifo2_writable;
assign hdmi2usbsoc_sdram_bankmachine2_syncfifo2_we = hdmi2usbsoc_sdram_bankmachine2_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine2_fifo_in_first = hdmi2usbsoc_sdram_bankmachine2_sink_first;
assign hdmi2usbsoc_sdram_bankmachine2_fifo_in_last = hdmi2usbsoc_sdram_bankmachine2_sink_last;
assign hdmi2usbsoc_sdram_bankmachine2_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine2_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine2_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine2_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine2_source_valid = hdmi2usbsoc_sdram_bankmachine2_syncfifo2_readable;
assign hdmi2usbsoc_sdram_bankmachine2_source_first = hdmi2usbsoc_sdram_bankmachine2_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine2_source_last = hdmi2usbsoc_sdram_bankmachine2_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine2_source_payload_we = hdmi2usbsoc_sdram_bankmachine2_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine2_source_payload_adr = hdmi2usbsoc_sdram_bankmachine2_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine2_syncfifo2_re = hdmi2usbsoc_sdram_bankmachine2_source_ready;

// synthesis translate_off
reg dummy_d_21;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine2_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine2_replace) begin
		hdmi2usbsoc_sdram_bankmachine2_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine2_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine2_wrport_adr <= hdmi2usbsoc_sdram_bankmachine2_produce;
	end
// synthesis translate_off
	dummy_d_21 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine2_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine2_syncfifo2_din;
assign hdmi2usbsoc_sdram_bankmachine2_wrport_we = (hdmi2usbsoc_sdram_bankmachine2_syncfifo2_we & (hdmi2usbsoc_sdram_bankmachine2_syncfifo2_writable | hdmi2usbsoc_sdram_bankmachine2_replace));
assign hdmi2usbsoc_sdram_bankmachine2_do_read = (hdmi2usbsoc_sdram_bankmachine2_syncfifo2_readable & hdmi2usbsoc_sdram_bankmachine2_syncfifo2_re);
assign hdmi2usbsoc_sdram_bankmachine2_rdport_adr = hdmi2usbsoc_sdram_bankmachine2_consume;
assign hdmi2usbsoc_sdram_bankmachine2_syncfifo2_dout = hdmi2usbsoc_sdram_bankmachine2_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine2_syncfifo2_writable = (hdmi2usbsoc_sdram_bankmachine2_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine2_syncfifo2_readable = (hdmi2usbsoc_sdram_bankmachine2_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine2_done = (hdmi2usbsoc_sdram_bankmachine2_count == 1'd0);

// synthesis translate_off
reg dummy_d_22;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine2_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_sel_row_adr <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_req_wdata_ready <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_req_rdata_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine2_cmd_valid <= 1'd0;
	controllerinjector_bankmachine2_next_state <= 3'd0;
	controllerinjector_bankmachine2_next_state <= controllerinjector_bankmachine2_state;
	case (controllerinjector_bankmachine2_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine2_done) begin
				hdmi2usbsoc_sdram_bankmachine2_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine2_cmd_ready) begin
					controllerinjector_bankmachine2_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine2_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine2_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine2_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine2_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine2_cmd_ready) begin
				controllerinjector_bankmachine2_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine2_done) begin
				hdmi2usbsoc_sdram_bankmachine2_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine2_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine2_refresh_req)) begin
				controllerinjector_bankmachine2_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine2_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine2_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine2_refresh_req) begin
				controllerinjector_bankmachine2_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine2_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine2_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine2_hit) begin
							hdmi2usbsoc_sdram_bankmachine2_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine2_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine2_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine2_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine2_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine2_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine2_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine2_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine2_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_22 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine3_sink_valid = hdmi2usbsoc_sdram_bankmachine3_req_valid;
assign hdmi2usbsoc_sdram_bankmachine3_req_ready = hdmi2usbsoc_sdram_bankmachine3_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine3_sink_payload_we = hdmi2usbsoc_sdram_bankmachine3_req_we;
assign hdmi2usbsoc_sdram_bankmachine3_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine3_req_adr;
assign hdmi2usbsoc_sdram_bankmachine3_source_ready = (hdmi2usbsoc_sdram_bankmachine3_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine3_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine3_req_lock = hdmi2usbsoc_sdram_bankmachine3_source_valid;
assign hdmi2usbsoc_sdram_bankmachine3_hit = (hdmi2usbsoc_sdram_bankmachine3_openrow == hdmi2usbsoc_sdram_bankmachine3_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ba = 2'd3;

// synthesis translate_off
reg dummy_d_23;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine3_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine3_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine3_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine3_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine3_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine3_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_23 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine3_wait = (~((hdmi2usbsoc_sdram_bankmachine3_cmd_valid & hdmi2usbsoc_sdram_bankmachine3_cmd_ready) & hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine3_syncfifo3_din = {hdmi2usbsoc_sdram_bankmachine3_fifo_in_last, hdmi2usbsoc_sdram_bankmachine3_fifo_in_first, hdmi2usbsoc_sdram_bankmachine3_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine3_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine3_fifo_out_last, hdmi2usbsoc_sdram_bankmachine3_fifo_out_first, hdmi2usbsoc_sdram_bankmachine3_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine3_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine3_syncfifo3_dout;
assign hdmi2usbsoc_sdram_bankmachine3_sink_ready = hdmi2usbsoc_sdram_bankmachine3_syncfifo3_writable;
assign hdmi2usbsoc_sdram_bankmachine3_syncfifo3_we = hdmi2usbsoc_sdram_bankmachine3_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine3_fifo_in_first = hdmi2usbsoc_sdram_bankmachine3_sink_first;
assign hdmi2usbsoc_sdram_bankmachine3_fifo_in_last = hdmi2usbsoc_sdram_bankmachine3_sink_last;
assign hdmi2usbsoc_sdram_bankmachine3_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine3_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine3_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine3_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine3_source_valid = hdmi2usbsoc_sdram_bankmachine3_syncfifo3_readable;
assign hdmi2usbsoc_sdram_bankmachine3_source_first = hdmi2usbsoc_sdram_bankmachine3_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine3_source_last = hdmi2usbsoc_sdram_bankmachine3_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine3_source_payload_we = hdmi2usbsoc_sdram_bankmachine3_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine3_source_payload_adr = hdmi2usbsoc_sdram_bankmachine3_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine3_syncfifo3_re = hdmi2usbsoc_sdram_bankmachine3_source_ready;

// synthesis translate_off
reg dummy_d_24;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine3_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine3_replace) begin
		hdmi2usbsoc_sdram_bankmachine3_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine3_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine3_wrport_adr <= hdmi2usbsoc_sdram_bankmachine3_produce;
	end
// synthesis translate_off
	dummy_d_24 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine3_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine3_syncfifo3_din;
assign hdmi2usbsoc_sdram_bankmachine3_wrport_we = (hdmi2usbsoc_sdram_bankmachine3_syncfifo3_we & (hdmi2usbsoc_sdram_bankmachine3_syncfifo3_writable | hdmi2usbsoc_sdram_bankmachine3_replace));
assign hdmi2usbsoc_sdram_bankmachine3_do_read = (hdmi2usbsoc_sdram_bankmachine3_syncfifo3_readable & hdmi2usbsoc_sdram_bankmachine3_syncfifo3_re);
assign hdmi2usbsoc_sdram_bankmachine3_rdport_adr = hdmi2usbsoc_sdram_bankmachine3_consume;
assign hdmi2usbsoc_sdram_bankmachine3_syncfifo3_dout = hdmi2usbsoc_sdram_bankmachine3_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine3_syncfifo3_writable = (hdmi2usbsoc_sdram_bankmachine3_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine3_syncfifo3_readable = (hdmi2usbsoc_sdram_bankmachine3_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine3_done = (hdmi2usbsoc_sdram_bankmachine3_count == 1'd0);

// synthesis translate_off
reg dummy_d_25;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine3_req_rdata_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_cmd_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ras <= 1'd0;
	controllerinjector_bankmachine3_next_state <= 3'd0;
	hdmi2usbsoc_sdram_bankmachine3_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_sel_row_adr <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine3_req_wdata_ready <= 1'd0;
	controllerinjector_bankmachine3_next_state <= controllerinjector_bankmachine3_state;
	case (controllerinjector_bankmachine3_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine3_done) begin
				hdmi2usbsoc_sdram_bankmachine3_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine3_cmd_ready) begin
					controllerinjector_bankmachine3_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine3_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine3_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine3_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine3_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine3_cmd_ready) begin
				controllerinjector_bankmachine3_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine3_done) begin
				hdmi2usbsoc_sdram_bankmachine3_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine3_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine3_refresh_req)) begin
				controllerinjector_bankmachine3_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine3_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine3_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine3_refresh_req) begin
				controllerinjector_bankmachine3_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine3_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine3_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine3_hit) begin
							hdmi2usbsoc_sdram_bankmachine3_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine3_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine3_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine3_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine3_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine3_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine3_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine3_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine3_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_25 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine4_sink_valid = hdmi2usbsoc_sdram_bankmachine4_req_valid;
assign hdmi2usbsoc_sdram_bankmachine4_req_ready = hdmi2usbsoc_sdram_bankmachine4_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine4_sink_payload_we = hdmi2usbsoc_sdram_bankmachine4_req_we;
assign hdmi2usbsoc_sdram_bankmachine4_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine4_req_adr;
assign hdmi2usbsoc_sdram_bankmachine4_source_ready = (hdmi2usbsoc_sdram_bankmachine4_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine4_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine4_req_lock = hdmi2usbsoc_sdram_bankmachine4_source_valid;
assign hdmi2usbsoc_sdram_bankmachine4_hit = (hdmi2usbsoc_sdram_bankmachine4_openrow == hdmi2usbsoc_sdram_bankmachine4_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ba = 3'd4;

// synthesis translate_off
reg dummy_d_26;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine4_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine4_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine4_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine4_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine4_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine4_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_26 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine4_wait = (~((hdmi2usbsoc_sdram_bankmachine4_cmd_valid & hdmi2usbsoc_sdram_bankmachine4_cmd_ready) & hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine4_syncfifo4_din = {hdmi2usbsoc_sdram_bankmachine4_fifo_in_last, hdmi2usbsoc_sdram_bankmachine4_fifo_in_first, hdmi2usbsoc_sdram_bankmachine4_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine4_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine4_fifo_out_last, hdmi2usbsoc_sdram_bankmachine4_fifo_out_first, hdmi2usbsoc_sdram_bankmachine4_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine4_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine4_syncfifo4_dout;
assign hdmi2usbsoc_sdram_bankmachine4_sink_ready = hdmi2usbsoc_sdram_bankmachine4_syncfifo4_writable;
assign hdmi2usbsoc_sdram_bankmachine4_syncfifo4_we = hdmi2usbsoc_sdram_bankmachine4_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine4_fifo_in_first = hdmi2usbsoc_sdram_bankmachine4_sink_first;
assign hdmi2usbsoc_sdram_bankmachine4_fifo_in_last = hdmi2usbsoc_sdram_bankmachine4_sink_last;
assign hdmi2usbsoc_sdram_bankmachine4_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine4_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine4_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine4_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine4_source_valid = hdmi2usbsoc_sdram_bankmachine4_syncfifo4_readable;
assign hdmi2usbsoc_sdram_bankmachine4_source_first = hdmi2usbsoc_sdram_bankmachine4_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine4_source_last = hdmi2usbsoc_sdram_bankmachine4_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine4_source_payload_we = hdmi2usbsoc_sdram_bankmachine4_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine4_source_payload_adr = hdmi2usbsoc_sdram_bankmachine4_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine4_syncfifo4_re = hdmi2usbsoc_sdram_bankmachine4_source_ready;

// synthesis translate_off
reg dummy_d_27;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine4_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine4_replace) begin
		hdmi2usbsoc_sdram_bankmachine4_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine4_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine4_wrport_adr <= hdmi2usbsoc_sdram_bankmachine4_produce;
	end
// synthesis translate_off
	dummy_d_27 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine4_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine4_syncfifo4_din;
assign hdmi2usbsoc_sdram_bankmachine4_wrport_we = (hdmi2usbsoc_sdram_bankmachine4_syncfifo4_we & (hdmi2usbsoc_sdram_bankmachine4_syncfifo4_writable | hdmi2usbsoc_sdram_bankmachine4_replace));
assign hdmi2usbsoc_sdram_bankmachine4_do_read = (hdmi2usbsoc_sdram_bankmachine4_syncfifo4_readable & hdmi2usbsoc_sdram_bankmachine4_syncfifo4_re);
assign hdmi2usbsoc_sdram_bankmachine4_rdport_adr = hdmi2usbsoc_sdram_bankmachine4_consume;
assign hdmi2usbsoc_sdram_bankmachine4_syncfifo4_dout = hdmi2usbsoc_sdram_bankmachine4_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine4_syncfifo4_writable = (hdmi2usbsoc_sdram_bankmachine4_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine4_syncfifo4_readable = (hdmi2usbsoc_sdram_bankmachine4_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine4_done = (hdmi2usbsoc_sdram_bankmachine4_count == 1'd0);

// synthesis translate_off
reg dummy_d_28;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine4_req_wdata_ready <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_req_rdata_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_cmd_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_sel_row_adr <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd0;
	controllerinjector_bankmachine4_next_state <= 3'd0;
	controllerinjector_bankmachine4_next_state <= controllerinjector_bankmachine4_state;
	case (controllerinjector_bankmachine4_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine4_done) begin
				hdmi2usbsoc_sdram_bankmachine4_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine4_cmd_ready) begin
					controllerinjector_bankmachine4_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine4_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine4_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine4_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine4_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine4_cmd_ready) begin
				controllerinjector_bankmachine4_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine4_done) begin
				hdmi2usbsoc_sdram_bankmachine4_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine4_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine4_refresh_req)) begin
				controllerinjector_bankmachine4_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine4_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine4_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine4_refresh_req) begin
				controllerinjector_bankmachine4_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine4_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine4_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine4_hit) begin
							hdmi2usbsoc_sdram_bankmachine4_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine4_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine4_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine4_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine4_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine4_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine4_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine4_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine4_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_28 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine5_sink_valid = hdmi2usbsoc_sdram_bankmachine5_req_valid;
assign hdmi2usbsoc_sdram_bankmachine5_req_ready = hdmi2usbsoc_sdram_bankmachine5_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine5_sink_payload_we = hdmi2usbsoc_sdram_bankmachine5_req_we;
assign hdmi2usbsoc_sdram_bankmachine5_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine5_req_adr;
assign hdmi2usbsoc_sdram_bankmachine5_source_ready = (hdmi2usbsoc_sdram_bankmachine5_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine5_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine5_req_lock = hdmi2usbsoc_sdram_bankmachine5_source_valid;
assign hdmi2usbsoc_sdram_bankmachine5_hit = (hdmi2usbsoc_sdram_bankmachine5_openrow == hdmi2usbsoc_sdram_bankmachine5_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ba = 3'd5;

// synthesis translate_off
reg dummy_d_29;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine5_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine5_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine5_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine5_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine5_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine5_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_29 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine5_wait = (~((hdmi2usbsoc_sdram_bankmachine5_cmd_valid & hdmi2usbsoc_sdram_bankmachine5_cmd_ready) & hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine5_syncfifo5_din = {hdmi2usbsoc_sdram_bankmachine5_fifo_in_last, hdmi2usbsoc_sdram_bankmachine5_fifo_in_first, hdmi2usbsoc_sdram_bankmachine5_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine5_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine5_fifo_out_last, hdmi2usbsoc_sdram_bankmachine5_fifo_out_first, hdmi2usbsoc_sdram_bankmachine5_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine5_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine5_syncfifo5_dout;
assign hdmi2usbsoc_sdram_bankmachine5_sink_ready = hdmi2usbsoc_sdram_bankmachine5_syncfifo5_writable;
assign hdmi2usbsoc_sdram_bankmachine5_syncfifo5_we = hdmi2usbsoc_sdram_bankmachine5_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine5_fifo_in_first = hdmi2usbsoc_sdram_bankmachine5_sink_first;
assign hdmi2usbsoc_sdram_bankmachine5_fifo_in_last = hdmi2usbsoc_sdram_bankmachine5_sink_last;
assign hdmi2usbsoc_sdram_bankmachine5_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine5_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine5_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine5_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine5_source_valid = hdmi2usbsoc_sdram_bankmachine5_syncfifo5_readable;
assign hdmi2usbsoc_sdram_bankmachine5_source_first = hdmi2usbsoc_sdram_bankmachine5_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine5_source_last = hdmi2usbsoc_sdram_bankmachine5_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine5_source_payload_we = hdmi2usbsoc_sdram_bankmachine5_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine5_source_payload_adr = hdmi2usbsoc_sdram_bankmachine5_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine5_syncfifo5_re = hdmi2usbsoc_sdram_bankmachine5_source_ready;

// synthesis translate_off
reg dummy_d_30;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine5_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine5_replace) begin
		hdmi2usbsoc_sdram_bankmachine5_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine5_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine5_wrport_adr <= hdmi2usbsoc_sdram_bankmachine5_produce;
	end
// synthesis translate_off
	dummy_d_30 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine5_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine5_syncfifo5_din;
assign hdmi2usbsoc_sdram_bankmachine5_wrport_we = (hdmi2usbsoc_sdram_bankmachine5_syncfifo5_we & (hdmi2usbsoc_sdram_bankmachine5_syncfifo5_writable | hdmi2usbsoc_sdram_bankmachine5_replace));
assign hdmi2usbsoc_sdram_bankmachine5_do_read = (hdmi2usbsoc_sdram_bankmachine5_syncfifo5_readable & hdmi2usbsoc_sdram_bankmachine5_syncfifo5_re);
assign hdmi2usbsoc_sdram_bankmachine5_rdport_adr = hdmi2usbsoc_sdram_bankmachine5_consume;
assign hdmi2usbsoc_sdram_bankmachine5_syncfifo5_dout = hdmi2usbsoc_sdram_bankmachine5_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine5_syncfifo5_writable = (hdmi2usbsoc_sdram_bankmachine5_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine5_syncfifo5_readable = (hdmi2usbsoc_sdram_bankmachine5_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine5_done = (hdmi2usbsoc_sdram_bankmachine5_count == 1'd0);

// synthesis translate_off
reg dummy_d_31;
// synthesis translate_on
always @(*) begin
	controllerinjector_bankmachine5_next_state <= 3'd0;
	hdmi2usbsoc_sdram_bankmachine5_req_wdata_ready <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_req_rdata_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_cmd_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_sel_row_adr <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd0;
	controllerinjector_bankmachine5_next_state <= controllerinjector_bankmachine5_state;
	case (controllerinjector_bankmachine5_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine5_done) begin
				hdmi2usbsoc_sdram_bankmachine5_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine5_cmd_ready) begin
					controllerinjector_bankmachine5_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine5_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine5_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine5_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine5_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine5_cmd_ready) begin
				controllerinjector_bankmachine5_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine5_done) begin
				hdmi2usbsoc_sdram_bankmachine5_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine5_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine5_refresh_req)) begin
				controllerinjector_bankmachine5_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine5_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine5_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine5_refresh_req) begin
				controllerinjector_bankmachine5_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine5_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine5_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine5_hit) begin
							hdmi2usbsoc_sdram_bankmachine5_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine5_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine5_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine5_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine5_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine5_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine5_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine5_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine5_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_31 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine6_sink_valid = hdmi2usbsoc_sdram_bankmachine6_req_valid;
assign hdmi2usbsoc_sdram_bankmachine6_req_ready = hdmi2usbsoc_sdram_bankmachine6_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine6_sink_payload_we = hdmi2usbsoc_sdram_bankmachine6_req_we;
assign hdmi2usbsoc_sdram_bankmachine6_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine6_req_adr;
assign hdmi2usbsoc_sdram_bankmachine6_source_ready = (hdmi2usbsoc_sdram_bankmachine6_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine6_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine6_req_lock = hdmi2usbsoc_sdram_bankmachine6_source_valid;
assign hdmi2usbsoc_sdram_bankmachine6_hit = (hdmi2usbsoc_sdram_bankmachine6_openrow == hdmi2usbsoc_sdram_bankmachine6_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ba = 3'd6;

// synthesis translate_off
reg dummy_d_32;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine6_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine6_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine6_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine6_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine6_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine6_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_32 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine6_wait = (~((hdmi2usbsoc_sdram_bankmachine6_cmd_valid & hdmi2usbsoc_sdram_bankmachine6_cmd_ready) & hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine6_syncfifo6_din = {hdmi2usbsoc_sdram_bankmachine6_fifo_in_last, hdmi2usbsoc_sdram_bankmachine6_fifo_in_first, hdmi2usbsoc_sdram_bankmachine6_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine6_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine6_fifo_out_last, hdmi2usbsoc_sdram_bankmachine6_fifo_out_first, hdmi2usbsoc_sdram_bankmachine6_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine6_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine6_syncfifo6_dout;
assign hdmi2usbsoc_sdram_bankmachine6_sink_ready = hdmi2usbsoc_sdram_bankmachine6_syncfifo6_writable;
assign hdmi2usbsoc_sdram_bankmachine6_syncfifo6_we = hdmi2usbsoc_sdram_bankmachine6_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine6_fifo_in_first = hdmi2usbsoc_sdram_bankmachine6_sink_first;
assign hdmi2usbsoc_sdram_bankmachine6_fifo_in_last = hdmi2usbsoc_sdram_bankmachine6_sink_last;
assign hdmi2usbsoc_sdram_bankmachine6_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine6_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine6_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine6_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine6_source_valid = hdmi2usbsoc_sdram_bankmachine6_syncfifo6_readable;
assign hdmi2usbsoc_sdram_bankmachine6_source_first = hdmi2usbsoc_sdram_bankmachine6_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine6_source_last = hdmi2usbsoc_sdram_bankmachine6_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine6_source_payload_we = hdmi2usbsoc_sdram_bankmachine6_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine6_source_payload_adr = hdmi2usbsoc_sdram_bankmachine6_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine6_syncfifo6_re = hdmi2usbsoc_sdram_bankmachine6_source_ready;

// synthesis translate_off
reg dummy_d_33;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine6_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine6_replace) begin
		hdmi2usbsoc_sdram_bankmachine6_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine6_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine6_wrport_adr <= hdmi2usbsoc_sdram_bankmachine6_produce;
	end
// synthesis translate_off
	dummy_d_33 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine6_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine6_syncfifo6_din;
assign hdmi2usbsoc_sdram_bankmachine6_wrport_we = (hdmi2usbsoc_sdram_bankmachine6_syncfifo6_we & (hdmi2usbsoc_sdram_bankmachine6_syncfifo6_writable | hdmi2usbsoc_sdram_bankmachine6_replace));
assign hdmi2usbsoc_sdram_bankmachine6_do_read = (hdmi2usbsoc_sdram_bankmachine6_syncfifo6_readable & hdmi2usbsoc_sdram_bankmachine6_syncfifo6_re);
assign hdmi2usbsoc_sdram_bankmachine6_rdport_adr = hdmi2usbsoc_sdram_bankmachine6_consume;
assign hdmi2usbsoc_sdram_bankmachine6_syncfifo6_dout = hdmi2usbsoc_sdram_bankmachine6_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine6_syncfifo6_writable = (hdmi2usbsoc_sdram_bankmachine6_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine6_syncfifo6_readable = (hdmi2usbsoc_sdram_bankmachine6_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine6_done = (hdmi2usbsoc_sdram_bankmachine6_count == 1'd0);

// synthesis translate_off
reg dummy_d_34;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd0;
	controllerinjector_bankmachine6_next_state <= 3'd0;
	hdmi2usbsoc_sdram_bankmachine6_req_wdata_ready <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_req_rdata_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_cmd_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_sel_row_adr <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd0;
	controllerinjector_bankmachine6_next_state <= controllerinjector_bankmachine6_state;
	case (controllerinjector_bankmachine6_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine6_done) begin
				hdmi2usbsoc_sdram_bankmachine6_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine6_cmd_ready) begin
					controllerinjector_bankmachine6_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine6_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine6_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine6_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine6_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine6_cmd_ready) begin
				controllerinjector_bankmachine6_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine6_done) begin
				hdmi2usbsoc_sdram_bankmachine6_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine6_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine6_refresh_req)) begin
				controllerinjector_bankmachine6_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine6_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine6_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine6_refresh_req) begin
				controllerinjector_bankmachine6_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine6_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine6_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine6_hit) begin
							hdmi2usbsoc_sdram_bankmachine6_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine6_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine6_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine6_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine6_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine6_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine6_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine6_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine6_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_34 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine7_sink_valid = hdmi2usbsoc_sdram_bankmachine7_req_valid;
assign hdmi2usbsoc_sdram_bankmachine7_req_ready = hdmi2usbsoc_sdram_bankmachine7_sink_ready;
assign hdmi2usbsoc_sdram_bankmachine7_sink_payload_we = hdmi2usbsoc_sdram_bankmachine7_req_we;
assign hdmi2usbsoc_sdram_bankmachine7_sink_payload_adr = hdmi2usbsoc_sdram_bankmachine7_req_adr;
assign hdmi2usbsoc_sdram_bankmachine7_source_ready = (hdmi2usbsoc_sdram_bankmachine7_req_wdata_ready | hdmi2usbsoc_sdram_bankmachine7_req_rdata_valid);
assign hdmi2usbsoc_sdram_bankmachine7_req_lock = hdmi2usbsoc_sdram_bankmachine7_source_valid;
assign hdmi2usbsoc_sdram_bankmachine7_hit = (hdmi2usbsoc_sdram_bankmachine7_openrow == hdmi2usbsoc_sdram_bankmachine7_source_payload_adr[20:8]);
assign hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ba = 3'd7;

// synthesis translate_off
reg dummy_d_35;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine7_cmd_payload_a <= 13'd0;
	if (hdmi2usbsoc_sdram_bankmachine7_sel_row_adr) begin
		hdmi2usbsoc_sdram_bankmachine7_cmd_payload_a <= hdmi2usbsoc_sdram_bankmachine7_source_payload_adr[20:8];
	end else begin
		hdmi2usbsoc_sdram_bankmachine7_cmd_payload_a <= {hdmi2usbsoc_sdram_bankmachine7_source_payload_adr[7:0], {2{1'd0}}};
	end
// synthesis translate_off
	dummy_d_35 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine7_wait = (~((hdmi2usbsoc_sdram_bankmachine7_cmd_valid & hdmi2usbsoc_sdram_bankmachine7_cmd_ready) & hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_bankmachine7_syncfifo7_din = {hdmi2usbsoc_sdram_bankmachine7_fifo_in_last, hdmi2usbsoc_sdram_bankmachine7_fifo_in_first, hdmi2usbsoc_sdram_bankmachine7_fifo_in_payload_adr, hdmi2usbsoc_sdram_bankmachine7_fifo_in_payload_we};
assign {hdmi2usbsoc_sdram_bankmachine7_fifo_out_last, hdmi2usbsoc_sdram_bankmachine7_fifo_out_first, hdmi2usbsoc_sdram_bankmachine7_fifo_out_payload_adr, hdmi2usbsoc_sdram_bankmachine7_fifo_out_payload_we} = hdmi2usbsoc_sdram_bankmachine7_syncfifo7_dout;
assign hdmi2usbsoc_sdram_bankmachine7_sink_ready = hdmi2usbsoc_sdram_bankmachine7_syncfifo7_writable;
assign hdmi2usbsoc_sdram_bankmachine7_syncfifo7_we = hdmi2usbsoc_sdram_bankmachine7_sink_valid;
assign hdmi2usbsoc_sdram_bankmachine7_fifo_in_first = hdmi2usbsoc_sdram_bankmachine7_sink_first;
assign hdmi2usbsoc_sdram_bankmachine7_fifo_in_last = hdmi2usbsoc_sdram_bankmachine7_sink_last;
assign hdmi2usbsoc_sdram_bankmachine7_fifo_in_payload_we = hdmi2usbsoc_sdram_bankmachine7_sink_payload_we;
assign hdmi2usbsoc_sdram_bankmachine7_fifo_in_payload_adr = hdmi2usbsoc_sdram_bankmachine7_sink_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine7_source_valid = hdmi2usbsoc_sdram_bankmachine7_syncfifo7_readable;
assign hdmi2usbsoc_sdram_bankmachine7_source_first = hdmi2usbsoc_sdram_bankmachine7_fifo_out_first;
assign hdmi2usbsoc_sdram_bankmachine7_source_last = hdmi2usbsoc_sdram_bankmachine7_fifo_out_last;
assign hdmi2usbsoc_sdram_bankmachine7_source_payload_we = hdmi2usbsoc_sdram_bankmachine7_fifo_out_payload_we;
assign hdmi2usbsoc_sdram_bankmachine7_source_payload_adr = hdmi2usbsoc_sdram_bankmachine7_fifo_out_payload_adr;
assign hdmi2usbsoc_sdram_bankmachine7_syncfifo7_re = hdmi2usbsoc_sdram_bankmachine7_source_ready;

// synthesis translate_off
reg dummy_d_36;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine7_wrport_adr <= 3'd0;
	if (hdmi2usbsoc_sdram_bankmachine7_replace) begin
		hdmi2usbsoc_sdram_bankmachine7_wrport_adr <= (hdmi2usbsoc_sdram_bankmachine7_produce - 1'd1);
	end else begin
		hdmi2usbsoc_sdram_bankmachine7_wrport_adr <= hdmi2usbsoc_sdram_bankmachine7_produce;
	end
// synthesis translate_off
	dummy_d_36 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_bankmachine7_wrport_dat_w = hdmi2usbsoc_sdram_bankmachine7_syncfifo7_din;
assign hdmi2usbsoc_sdram_bankmachine7_wrport_we = (hdmi2usbsoc_sdram_bankmachine7_syncfifo7_we & (hdmi2usbsoc_sdram_bankmachine7_syncfifo7_writable | hdmi2usbsoc_sdram_bankmachine7_replace));
assign hdmi2usbsoc_sdram_bankmachine7_do_read = (hdmi2usbsoc_sdram_bankmachine7_syncfifo7_readable & hdmi2usbsoc_sdram_bankmachine7_syncfifo7_re);
assign hdmi2usbsoc_sdram_bankmachine7_rdport_adr = hdmi2usbsoc_sdram_bankmachine7_consume;
assign hdmi2usbsoc_sdram_bankmachine7_syncfifo7_dout = hdmi2usbsoc_sdram_bankmachine7_rdport_dat_r;
assign hdmi2usbsoc_sdram_bankmachine7_syncfifo7_writable = (hdmi2usbsoc_sdram_bankmachine7_level != 4'd8);
assign hdmi2usbsoc_sdram_bankmachine7_syncfifo7_readable = (hdmi2usbsoc_sdram_bankmachine7_level != 1'd0);
assign hdmi2usbsoc_sdram_bankmachine7_done = (hdmi2usbsoc_sdram_bankmachine7_count == 1'd0);

// synthesis translate_off
reg dummy_d_37;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine7_track_open <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_track_close <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_sel_row_adr <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd0;
	controllerinjector_bankmachine7_next_state <= 3'd0;
	hdmi2usbsoc_sdram_bankmachine7_req_wdata_ready <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_req_rdata_valid <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_refresh_gnt <= 1'd0;
	hdmi2usbsoc_sdram_bankmachine7_cmd_valid <= 1'd0;
	controllerinjector_bankmachine7_next_state <= controllerinjector_bankmachine7_state;
	case (controllerinjector_bankmachine7_state)
		1'd1: begin
			if (hdmi2usbsoc_sdram_bankmachine7_done) begin
				hdmi2usbsoc_sdram_bankmachine7_cmd_valid <= 1'd1;
				if (hdmi2usbsoc_sdram_bankmachine7_cmd_ready) begin
					controllerinjector_bankmachine7_next_state <= 3'd4;
				end
				hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
				hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine7_track_close <= 1'd1;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_bankmachine7_sel_row_adr <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine7_track_open <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine7_cmd_valid <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if (hdmi2usbsoc_sdram_bankmachine7_cmd_ready) begin
				controllerinjector_bankmachine7_next_state <= 3'd5;
			end
			hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (hdmi2usbsoc_sdram_bankmachine7_done) begin
				hdmi2usbsoc_sdram_bankmachine7_refresh_gnt <= 1'd1;
			end
			hdmi2usbsoc_sdram_bankmachine7_track_close <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if ((~hdmi2usbsoc_sdram_bankmachine7_refresh_req)) begin
				controllerinjector_bankmachine7_next_state <= 1'd0;
			end
		end
		3'd4: begin
			controllerinjector_bankmachine7_next_state <= 2'd2;
		end
		3'd5: begin
			controllerinjector_bankmachine7_next_state <= 1'd0;
		end
		default: begin
			if (hdmi2usbsoc_sdram_bankmachine7_refresh_req) begin
				controllerinjector_bankmachine7_next_state <= 2'd3;
			end else begin
				if (hdmi2usbsoc_sdram_bankmachine7_source_valid) begin
					if (hdmi2usbsoc_sdram_bankmachine7_has_openrow) begin
						if (hdmi2usbsoc_sdram_bankmachine7_hit) begin
							hdmi2usbsoc_sdram_bankmachine7_cmd_valid <= 1'd1;
							if (hdmi2usbsoc_sdram_bankmachine7_source_payload_we) begin
								hdmi2usbsoc_sdram_bankmachine7_req_wdata_ready <= hdmi2usbsoc_sdram_bankmachine7_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd1;
								hdmi2usbsoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
							end else begin
								hdmi2usbsoc_sdram_bankmachine7_req_rdata_valid <= hdmi2usbsoc_sdram_bankmachine7_cmd_ready;
								hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd1;
							end
							hdmi2usbsoc_sdram_bankmachine7_cmd_payload_cas <= 1'd1;
						end else begin
							controllerinjector_bankmachine7_next_state <= 1'd1;
						end
					end else begin
						controllerinjector_bankmachine7_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_37 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_read_available = ((((((((hdmi2usbsoc_sdram_bankmachine0_cmd_valid & hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read) | (hdmi2usbsoc_sdram_bankmachine1_cmd_valid & hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read)) | (hdmi2usbsoc_sdram_bankmachine2_cmd_valid & hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read)) | (hdmi2usbsoc_sdram_bankmachine3_cmd_valid & hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read)) | (hdmi2usbsoc_sdram_bankmachine4_cmd_valid & hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read)) | (hdmi2usbsoc_sdram_bankmachine5_cmd_valid & hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read)) | (hdmi2usbsoc_sdram_bankmachine6_cmd_valid & hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read)) | (hdmi2usbsoc_sdram_bankmachine7_cmd_valid & hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read));
assign hdmi2usbsoc_sdram_write_available = ((((((((hdmi2usbsoc_sdram_bankmachine0_cmd_valid & hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write) | (hdmi2usbsoc_sdram_bankmachine1_cmd_valid & hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write)) | (hdmi2usbsoc_sdram_bankmachine2_cmd_valid & hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write)) | (hdmi2usbsoc_sdram_bankmachine3_cmd_valid & hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write)) | (hdmi2usbsoc_sdram_bankmachine4_cmd_valid & hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write)) | (hdmi2usbsoc_sdram_bankmachine5_cmd_valid & hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write)) | (hdmi2usbsoc_sdram_bankmachine6_cmd_valid & hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write)) | (hdmi2usbsoc_sdram_bankmachine7_cmd_valid & hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write));
assign hdmi2usbsoc_sdram_max_time0 = (hdmi2usbsoc_sdram_time0 == 1'd0);
assign hdmi2usbsoc_sdram_max_time1 = (hdmi2usbsoc_sdram_time1 == 1'd0);
assign hdmi2usbsoc_sdram_bankmachine0_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_bankmachine1_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_bankmachine2_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_bankmachine3_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_bankmachine4_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_bankmachine5_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_bankmachine6_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_bankmachine7_refresh_req = hdmi2usbsoc_sdram_cmd_valid;
assign hdmi2usbsoc_sdram_go_to_refresh = (((((((hdmi2usbsoc_sdram_bankmachine0_refresh_gnt & hdmi2usbsoc_sdram_bankmachine1_refresh_gnt) & hdmi2usbsoc_sdram_bankmachine2_refresh_gnt) & hdmi2usbsoc_sdram_bankmachine3_refresh_gnt) & hdmi2usbsoc_sdram_bankmachine4_refresh_gnt) & hdmi2usbsoc_sdram_bankmachine5_refresh_gnt) & hdmi2usbsoc_sdram_bankmachine6_refresh_gnt) & hdmi2usbsoc_sdram_bankmachine7_refresh_gnt);
assign hdmi2usbsoc_sdram_interface_rdata = {hdmi2usbsoc_sdram_dfi_p1_rddata, hdmi2usbsoc_sdram_dfi_p0_rddata};
assign {hdmi2usbsoc_sdram_dfi_p1_wrdata, hdmi2usbsoc_sdram_dfi_p0_wrdata} = hdmi2usbsoc_sdram_interface_wdata;
assign {hdmi2usbsoc_sdram_dfi_p1_wrdata_mask, hdmi2usbsoc_sdram_dfi_p0_wrdata_mask} = (~hdmi2usbsoc_sdram_interface_wdata_we);

// synthesis translate_off
reg dummy_d_38;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_cmd_valids <= 8'd0;
	hdmi2usbsoc_sdram_choose_cmd_valids[0] <= (hdmi2usbsoc_sdram_bankmachine0_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
	hdmi2usbsoc_sdram_choose_cmd_valids[1] <= (hdmi2usbsoc_sdram_bankmachine1_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
	hdmi2usbsoc_sdram_choose_cmd_valids[2] <= (hdmi2usbsoc_sdram_bankmachine2_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
	hdmi2usbsoc_sdram_choose_cmd_valids[3] <= (hdmi2usbsoc_sdram_bankmachine3_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
	hdmi2usbsoc_sdram_choose_cmd_valids[4] <= (hdmi2usbsoc_sdram_bankmachine4_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
	hdmi2usbsoc_sdram_choose_cmd_valids[5] <= (hdmi2usbsoc_sdram_bankmachine5_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
	hdmi2usbsoc_sdram_choose_cmd_valids[6] <= (hdmi2usbsoc_sdram_bankmachine6_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
	hdmi2usbsoc_sdram_choose_cmd_valids[7] <= (hdmi2usbsoc_sdram_bankmachine7_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_cmd_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_cmd_want_reads) & (hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_cmd_want_writes))));
// synthesis translate_off
	dummy_d_38 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_choose_cmd_request = hdmi2usbsoc_sdram_choose_cmd_valids;
assign hdmi2usbsoc_sdram_choose_cmd_cmd_valid = comb_rhs_array_muxed0;
assign hdmi2usbsoc_sdram_choose_cmd_cmd_payload_a = comb_rhs_array_muxed1;
assign hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ba = comb_rhs_array_muxed2;
assign hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_read = comb_rhs_array_muxed3;
assign hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_write = comb_rhs_array_muxed4;
assign hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_cmd = comb_rhs_array_muxed5;

// synthesis translate_off
reg dummy_d_39;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_cmd_cmd_payload_cas <= 1'd0;
	if (hdmi2usbsoc_sdram_choose_cmd_cmd_valid) begin
		hdmi2usbsoc_sdram_choose_cmd_cmd_payload_cas <= comb_t_array_muxed0;
	end
// synthesis translate_off
	dummy_d_39 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_40;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ras <= 1'd0;
	if (hdmi2usbsoc_sdram_choose_cmd_cmd_valid) begin
		hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ras <= comb_t_array_muxed1;
	end
// synthesis translate_off
	dummy_d_40 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_41;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_cmd_cmd_payload_we <= 1'd0;
	if (hdmi2usbsoc_sdram_choose_cmd_cmd_valid) begin
		hdmi2usbsoc_sdram_choose_cmd_cmd_payload_we <= comb_t_array_muxed2;
	end
// synthesis translate_off
	dummy_d_41 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_choose_cmd_ce = hdmi2usbsoc_sdram_choose_cmd_cmd_ready;

// synthesis translate_off
reg dummy_d_42;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_req_valids <= 8'd0;
	hdmi2usbsoc_sdram_choose_req_valids[0] <= (hdmi2usbsoc_sdram_bankmachine0_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
	hdmi2usbsoc_sdram_choose_req_valids[1] <= (hdmi2usbsoc_sdram_bankmachine1_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
	hdmi2usbsoc_sdram_choose_req_valids[2] <= (hdmi2usbsoc_sdram_bankmachine2_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
	hdmi2usbsoc_sdram_choose_req_valids[3] <= (hdmi2usbsoc_sdram_bankmachine3_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
	hdmi2usbsoc_sdram_choose_req_valids[4] <= (hdmi2usbsoc_sdram_bankmachine4_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
	hdmi2usbsoc_sdram_choose_req_valids[5] <= (hdmi2usbsoc_sdram_bankmachine5_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
	hdmi2usbsoc_sdram_choose_req_valids[6] <= (hdmi2usbsoc_sdram_bankmachine6_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
	hdmi2usbsoc_sdram_choose_req_valids[7] <= (hdmi2usbsoc_sdram_bankmachine7_cmd_valid & ((hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd & hdmi2usbsoc_sdram_choose_req_want_cmds) | ((hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read == hdmi2usbsoc_sdram_choose_req_want_reads) & (hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write == hdmi2usbsoc_sdram_choose_req_want_writes))));
// synthesis translate_off
	dummy_d_42 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_choose_req_request = hdmi2usbsoc_sdram_choose_req_valids;
assign hdmi2usbsoc_sdram_choose_req_cmd_valid = comb_rhs_array_muxed6;
assign hdmi2usbsoc_sdram_choose_req_cmd_payload_a = comb_rhs_array_muxed7;
assign hdmi2usbsoc_sdram_choose_req_cmd_payload_ba = comb_rhs_array_muxed8;
assign hdmi2usbsoc_sdram_choose_req_cmd_payload_is_read = comb_rhs_array_muxed9;
assign hdmi2usbsoc_sdram_choose_req_cmd_payload_is_write = comb_rhs_array_muxed10;
assign hdmi2usbsoc_sdram_choose_req_cmd_payload_is_cmd = comb_rhs_array_muxed11;

// synthesis translate_off
reg dummy_d_43;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_req_cmd_payload_cas <= 1'd0;
	if (hdmi2usbsoc_sdram_choose_req_cmd_valid) begin
		hdmi2usbsoc_sdram_choose_req_cmd_payload_cas <= comb_t_array_muxed3;
	end
// synthesis translate_off
	dummy_d_43 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_44;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_req_cmd_payload_ras <= 1'd0;
	if (hdmi2usbsoc_sdram_choose_req_cmd_valid) begin
		hdmi2usbsoc_sdram_choose_req_cmd_payload_ras <= comb_t_array_muxed4;
	end
// synthesis translate_off
	dummy_d_44 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_45;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_req_cmd_payload_we <= 1'd0;
	if (hdmi2usbsoc_sdram_choose_req_cmd_valid) begin
		hdmi2usbsoc_sdram_choose_req_cmd_payload_we <= comb_t_array_muxed5;
	end
// synthesis translate_off
	dummy_d_45 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_46;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine0_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 1'd0))) begin
		hdmi2usbsoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 1'd0))) begin
		hdmi2usbsoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_46 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_47;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine1_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 1'd1))) begin
		hdmi2usbsoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 1'd1))) begin
		hdmi2usbsoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_47 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_48;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine2_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 2'd2))) begin
		hdmi2usbsoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 2'd2))) begin
		hdmi2usbsoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_48 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_49;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine3_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 2'd3))) begin
		hdmi2usbsoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 2'd3))) begin
		hdmi2usbsoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_49 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_50;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine4_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 3'd4))) begin
		hdmi2usbsoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 3'd4))) begin
		hdmi2usbsoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_50 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_51;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine5_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 3'd5))) begin
		hdmi2usbsoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 3'd5))) begin
		hdmi2usbsoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_51 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_52;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine6_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 3'd6))) begin
		hdmi2usbsoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 3'd6))) begin
		hdmi2usbsoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_52 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_53;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_bankmachine7_cmd_ready <= 1'd0;
	if (((hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_ready) & (hdmi2usbsoc_sdram_choose_cmd_grant == 3'd7))) begin
		hdmi2usbsoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
	if (((hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_ready) & (hdmi2usbsoc_sdram_choose_req_grant == 3'd7))) begin
		hdmi2usbsoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
// synthesis translate_off
	dummy_d_53 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sdram_choose_req_ce = hdmi2usbsoc_sdram_choose_req_cmd_ready;
assign hdmi2usbsoc_sdram_dfi_p0_cke = 1'd1;
assign hdmi2usbsoc_sdram_dfi_p0_cs_n = 1'd0;
assign hdmi2usbsoc_sdram_dfi_p0_odt = 1'd1;
assign hdmi2usbsoc_sdram_dfi_p0_reset_n = 1'd1;
assign hdmi2usbsoc_sdram_dfi_p1_cke = 1'd1;
assign hdmi2usbsoc_sdram_dfi_p1_cs_n = 1'd0;
assign hdmi2usbsoc_sdram_dfi_p1_odt = 1'd1;
assign hdmi2usbsoc_sdram_dfi_p1_reset_n = 1'd1;

// synthesis translate_off
reg dummy_d_54;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_choose_req_want_writes <= 1'd0;
	controllerinjector_multiplexer_next_state <= 4'd0;
	hdmi2usbsoc_sdram_choose_req_cmd_ready <= 1'd0;
	hdmi2usbsoc_sdram_cmd_ready <= 1'd0;
	hdmi2usbsoc_sdram_sel0 <= 2'd0;
	hdmi2usbsoc_sdram_sel1 <= 2'd0;
	hdmi2usbsoc_sdram_en0 <= 1'd0;
	hdmi2usbsoc_sdram_en1 <= 1'd0;
	hdmi2usbsoc_sdram_choose_cmd_cmd_ready <= 1'd0;
	hdmi2usbsoc_sdram_choose_req_want_reads <= 1'd0;
	controllerinjector_multiplexer_next_state <= controllerinjector_multiplexer_state;
	case (controllerinjector_multiplexer_state)
		1'd1: begin
			hdmi2usbsoc_sdram_en1 <= 1'd1;
			hdmi2usbsoc_sdram_choose_req_want_writes <= 1'd1;
			hdmi2usbsoc_sdram_choose_cmd_cmd_ready <= 1'd1;
			hdmi2usbsoc_sdram_choose_req_cmd_ready <= 1'd1;
			hdmi2usbsoc_sdram_sel0 <= 1'd1;
			hdmi2usbsoc_sdram_sel1 <= 2'd2;
			if (hdmi2usbsoc_sdram_read_available) begin
				if (((~hdmi2usbsoc_sdram_write_available) | hdmi2usbsoc_sdram_max_time1)) begin
					controllerinjector_multiplexer_next_state <= 3'd7;
				end
			end
			if (hdmi2usbsoc_sdram_go_to_refresh) begin
				controllerinjector_multiplexer_next_state <= 2'd2;
			end
		end
		2'd2: begin
			hdmi2usbsoc_sdram_sel0 <= 2'd3;
			hdmi2usbsoc_sdram_cmd_ready <= 1'd1;
			if (hdmi2usbsoc_sdram_cmd_last) begin
				controllerinjector_multiplexer_next_state <= 1'd0;
			end
		end
		2'd3: begin
			controllerinjector_multiplexer_next_state <= 3'd4;
		end
		3'd4: begin
			controllerinjector_multiplexer_next_state <= 3'd5;
		end
		3'd5: begin
			controllerinjector_multiplexer_next_state <= 3'd6;
		end
		3'd6: begin
			controllerinjector_multiplexer_next_state <= 1'd1;
		end
		3'd7: begin
			controllerinjector_multiplexer_next_state <= 4'd8;
		end
		4'd8: begin
			controllerinjector_multiplexer_next_state <= 1'd0;
		end
		default: begin
			hdmi2usbsoc_sdram_en0 <= 1'd1;
			hdmi2usbsoc_sdram_choose_req_want_reads <= 1'd1;
			hdmi2usbsoc_sdram_choose_cmd_cmd_ready <= 1'd1;
			hdmi2usbsoc_sdram_choose_req_cmd_ready <= 1'd1;
			hdmi2usbsoc_sdram_sel0 <= 2'd2;
			hdmi2usbsoc_sdram_sel1 <= 1'd1;
			if (hdmi2usbsoc_sdram_write_available) begin
				if (((~hdmi2usbsoc_sdram_read_available) | hdmi2usbsoc_sdram_max_time0)) begin
					controllerinjector_multiplexer_next_state <= 2'd3;
				end
			end
			if (hdmi2usbsoc_sdram_go_to_refresh) begin
				controllerinjector_multiplexer_next_state <= 2'd2;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_54 <= dummy_s;
// synthesis translate_on
end
assign controllerinjector_cba0 = hdmi2usbsoc_port_cmd_payload_adr[10:8];
assign controllerinjector_rca0 = {hdmi2usbsoc_port_cmd_payload_adr[23:11], hdmi2usbsoc_port_cmd_payload_adr[7:0]};
assign controllerinjector_cba1 = hdmi2usbsoc_litedramport0_cmd_payload_adr0[10:8];
assign controllerinjector_rca1 = {hdmi2usbsoc_litedramport0_cmd_payload_adr0[23:11], hdmi2usbsoc_litedramport0_cmd_payload_adr0[7:0]};
assign controllerinjector_cba2 = hdmi2usbsoc_litedramport1_cmd_payload_adr0[10:8];
assign controllerinjector_rca2 = {hdmi2usbsoc_litedramport1_cmd_payload_adr0[23:11], hdmi2usbsoc_litedramport1_cmd_payload_adr0[7:0]};
assign controllerinjector_cba3 = hdmi2usbsoc_litedramport2_cmd_payload_adr0[10:8];
assign controllerinjector_rca3 = {hdmi2usbsoc_litedramport2_cmd_payload_adr0[23:11], hdmi2usbsoc_litedramport2_cmd_payload_adr0[7:0]};
assign controllerinjector_cba4 = hdmi2usbsoc_litedramport3_cmd_payload_adr0[10:8];
assign controllerinjector_rca4 = {hdmi2usbsoc_litedramport3_cmd_payload_adr0[23:11], hdmi2usbsoc_litedramport3_cmd_payload_adr0[7:0]};
assign controllerinjector_cba5 = encoder_port_port_cmd_payload_adr[10:8];
assign controllerinjector_rca5 = {encoder_port_port_cmd_payload_adr[23:11], encoder_port_port_cmd_payload_adr[7:0]};
assign controllerinjector_roundrobin0_request = {(((controllerinjector_cba5 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin0_ce = ((~hdmi2usbsoc_sdram_interface_bank0_valid) & (~hdmi2usbsoc_sdram_interface_bank0_lock));
assign hdmi2usbsoc_sdram_interface_bank0_adr = comb_rhs_array_muxed12;
assign hdmi2usbsoc_sdram_interface_bank0_we = comb_rhs_array_muxed13;
assign hdmi2usbsoc_sdram_interface_bank0_valid = comb_rhs_array_muxed14;
assign controllerinjector_roundrobin1_request = {(((controllerinjector_cba5 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin1_ce = ((~hdmi2usbsoc_sdram_interface_bank1_valid) & (~hdmi2usbsoc_sdram_interface_bank1_lock));
assign hdmi2usbsoc_sdram_interface_bank1_adr = comb_rhs_array_muxed15;
assign hdmi2usbsoc_sdram_interface_bank1_we = comb_rhs_array_muxed16;
assign hdmi2usbsoc_sdram_interface_bank1_valid = comb_rhs_array_muxed17;
assign controllerinjector_roundrobin2_request = {(((controllerinjector_cba5 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin2_ce = ((~hdmi2usbsoc_sdram_interface_bank2_valid) & (~hdmi2usbsoc_sdram_interface_bank2_lock));
assign hdmi2usbsoc_sdram_interface_bank2_adr = comb_rhs_array_muxed18;
assign hdmi2usbsoc_sdram_interface_bank2_we = comb_rhs_array_muxed19;
assign hdmi2usbsoc_sdram_interface_bank2_valid = comb_rhs_array_muxed20;
assign controllerinjector_roundrobin3_request = {(((controllerinjector_cba5 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin3_ce = ((~hdmi2usbsoc_sdram_interface_bank3_valid) & (~hdmi2usbsoc_sdram_interface_bank3_lock));
assign hdmi2usbsoc_sdram_interface_bank3_adr = comb_rhs_array_muxed21;
assign hdmi2usbsoc_sdram_interface_bank3_we = comb_rhs_array_muxed22;
assign hdmi2usbsoc_sdram_interface_bank3_valid = comb_rhs_array_muxed23;
assign controllerinjector_roundrobin4_request = {(((controllerinjector_cba5 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin4_ce = ((~hdmi2usbsoc_sdram_interface_bank4_valid) & (~hdmi2usbsoc_sdram_interface_bank4_lock));
assign hdmi2usbsoc_sdram_interface_bank4_adr = comb_rhs_array_muxed24;
assign hdmi2usbsoc_sdram_interface_bank4_we = comb_rhs_array_muxed25;
assign hdmi2usbsoc_sdram_interface_bank4_valid = comb_rhs_array_muxed26;
assign controllerinjector_roundrobin5_request = {(((controllerinjector_cba5 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin5_ce = ((~hdmi2usbsoc_sdram_interface_bank5_valid) & (~hdmi2usbsoc_sdram_interface_bank5_lock));
assign hdmi2usbsoc_sdram_interface_bank5_adr = comb_rhs_array_muxed27;
assign hdmi2usbsoc_sdram_interface_bank5_we = comb_rhs_array_muxed28;
assign hdmi2usbsoc_sdram_interface_bank5_valid = comb_rhs_array_muxed29;
assign controllerinjector_roundrobin6_request = {(((controllerinjector_cba5 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin6_ce = ((~hdmi2usbsoc_sdram_interface_bank6_valid) & (~hdmi2usbsoc_sdram_interface_bank6_lock));
assign hdmi2usbsoc_sdram_interface_bank6_adr = comb_rhs_array_muxed30;
assign hdmi2usbsoc_sdram_interface_bank6_we = comb_rhs_array_muxed31;
assign hdmi2usbsoc_sdram_interface_bank6_valid = comb_rhs_array_muxed32;
assign controllerinjector_roundrobin7_request = {(((controllerinjector_cba5 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))))) & encoder_port_port_cmd_valid), (((controllerinjector_cba4 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0), (((controllerinjector_cba3 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0), (((controllerinjector_cba2 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0), (((controllerinjector_cba1 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0), (((controllerinjector_cba0 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid)};
assign controllerinjector_roundrobin7_ce = ((~hdmi2usbsoc_sdram_interface_bank7_valid) & (~hdmi2usbsoc_sdram_interface_bank7_lock));
assign hdmi2usbsoc_sdram_interface_bank7_adr = comb_rhs_array_muxed33;
assign hdmi2usbsoc_sdram_interface_bank7_we = comb_rhs_array_muxed34;
assign hdmi2usbsoc_sdram_interface_bank7_valid = comb_rhs_array_muxed35;
assign hdmi2usbsoc_port_cmd_ready = ((((((((1'd0 | (((controllerinjector_roundrobin0_grant == 1'd0) & ((controllerinjector_cba0 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank0_ready)) | (((controllerinjector_roundrobin1_grant == 1'd0) & ((controllerinjector_cba0 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank1_ready)) | (((controllerinjector_roundrobin2_grant == 1'd0) & ((controllerinjector_cba0 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank2_ready)) | (((controllerinjector_roundrobin3_grant == 1'd0) & ((controllerinjector_cba0 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank3_ready)) | (((controllerinjector_roundrobin4_grant == 1'd0) & ((controllerinjector_cba0 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank4_ready)) | (((controllerinjector_roundrobin5_grant == 1'd0) & ((controllerinjector_cba0 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank5_ready)) | (((controllerinjector_roundrobin6_grant == 1'd0) & ((controllerinjector_cba0 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank6_ready)) | (((controllerinjector_roundrobin7_grant == 1'd0) & ((controllerinjector_cba0 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0)))))) & hdmi2usbsoc_sdram_interface_bank7_ready));
assign hdmi2usbsoc_litedramport0_cmd_ready0 = ((((((((1'd0 | (((controllerinjector_roundrobin0_grant == 1'd1) & ((controllerinjector_cba1 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank0_ready)) | (((controllerinjector_roundrobin1_grant == 1'd1) & ((controllerinjector_cba1 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank1_ready)) | (((controllerinjector_roundrobin2_grant == 1'd1) & ((controllerinjector_cba1 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank2_ready)) | (((controllerinjector_roundrobin3_grant == 1'd1) & ((controllerinjector_cba1 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank3_ready)) | (((controllerinjector_roundrobin4_grant == 1'd1) & ((controllerinjector_cba1 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank4_ready)) | (((controllerinjector_roundrobin5_grant == 1'd1) & ((controllerinjector_cba1 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank5_ready)) | (((controllerinjector_roundrobin6_grant == 1'd1) & ((controllerinjector_cba1 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank6_ready)) | (((controllerinjector_roundrobin7_grant == 1'd1) & ((controllerinjector_cba1 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1)))))) & hdmi2usbsoc_sdram_interface_bank7_ready));
assign hdmi2usbsoc_litedramport1_cmd_ready0 = ((((((((1'd0 | (((controllerinjector_roundrobin0_grant == 2'd2) & ((controllerinjector_cba2 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank0_ready)) | (((controllerinjector_roundrobin1_grant == 2'd2) & ((controllerinjector_cba2 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank1_ready)) | (((controllerinjector_roundrobin2_grant == 2'd2) & ((controllerinjector_cba2 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank2_ready)) | (((controllerinjector_roundrobin3_grant == 2'd2) & ((controllerinjector_cba2 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank3_ready)) | (((controllerinjector_roundrobin4_grant == 2'd2) & ((controllerinjector_cba2 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank4_ready)) | (((controllerinjector_roundrobin5_grant == 2'd2) & ((controllerinjector_cba2 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank5_ready)) | (((controllerinjector_roundrobin6_grant == 2'd2) & ((controllerinjector_cba2 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank6_ready)) | (((controllerinjector_roundrobin7_grant == 2'd2) & ((controllerinjector_cba2 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2)))))) & hdmi2usbsoc_sdram_interface_bank7_ready));
assign hdmi2usbsoc_litedramport2_cmd_ready0 = ((((((((1'd0 | (((controllerinjector_roundrobin0_grant == 2'd3) & ((controllerinjector_cba3 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank0_ready)) | (((controllerinjector_roundrobin1_grant == 2'd3) & ((controllerinjector_cba3 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank1_ready)) | (((controllerinjector_roundrobin2_grant == 2'd3) & ((controllerinjector_cba3 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank2_ready)) | (((controllerinjector_roundrobin3_grant == 2'd3) & ((controllerinjector_cba3 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank3_ready)) | (((controllerinjector_roundrobin4_grant == 2'd3) & ((controllerinjector_cba3 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank4_ready)) | (((controllerinjector_roundrobin5_grant == 2'd3) & ((controllerinjector_cba3 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank5_ready)) | (((controllerinjector_roundrobin6_grant == 2'd3) & ((controllerinjector_cba3 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank6_ready)) | (((controllerinjector_roundrobin7_grant == 2'd3) & ((controllerinjector_cba3 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3)))))) & hdmi2usbsoc_sdram_interface_bank7_ready));
assign hdmi2usbsoc_litedramport3_cmd_ready0 = ((((((((1'd0 | (((controllerinjector_roundrobin0_grant == 3'd4) & ((controllerinjector_cba4 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank0_ready)) | (((controllerinjector_roundrobin1_grant == 3'd4) & ((controllerinjector_cba4 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank1_ready)) | (((controllerinjector_roundrobin2_grant == 3'd4) & ((controllerinjector_cba4 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank2_ready)) | (((controllerinjector_roundrobin3_grant == 3'd4) & ((controllerinjector_cba4 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank3_ready)) | (((controllerinjector_roundrobin4_grant == 3'd4) & ((controllerinjector_cba4 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank4_ready)) | (((controllerinjector_roundrobin5_grant == 3'd4) & ((controllerinjector_cba4 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank5_ready)) | (((controllerinjector_roundrobin6_grant == 3'd4) & ((controllerinjector_cba4 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank6_ready)) | (((controllerinjector_roundrobin7_grant == 3'd4) & ((controllerinjector_cba4 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4)))))) & hdmi2usbsoc_sdram_interface_bank7_ready));
assign encoder_port_port_cmd_ready = ((((((((1'd0 | (((controllerinjector_roundrobin0_grant == 3'd5) & ((controllerinjector_cba5 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank0_ready)) | (((controllerinjector_roundrobin1_grant == 3'd5) & ((controllerinjector_cba5 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank1_ready)) | (((controllerinjector_roundrobin2_grant == 3'd5) & ((controllerinjector_cba5 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank2_ready)) | (((controllerinjector_roundrobin3_grant == 3'd5) & ((controllerinjector_cba5 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank3_ready)) | (((controllerinjector_roundrobin4_grant == 3'd5) & ((controllerinjector_cba5 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank4_ready)) | (((controllerinjector_roundrobin5_grant == 3'd5) & ((controllerinjector_cba5 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank5_ready)) | (((controllerinjector_roundrobin6_grant == 3'd5) & ((controllerinjector_cba5 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank6_ready)) | (((controllerinjector_roundrobin7_grant == 3'd5) & ((controllerinjector_cba5 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5)))))) & hdmi2usbsoc_sdram_interface_bank7_ready));
assign hdmi2usbsoc_port_wdata_ready = controllerinjector_new_master_wdata_ready0;
assign hdmi2usbsoc_litedramport0_wdata_ready = controllerinjector_new_master_wdata_ready1;
assign hdmi2usbsoc_litedramport1_wdata_ready = controllerinjector_new_master_wdata_ready2;
assign hdmi2usbsoc_litedramport2_wdata_ready = controllerinjector_new_master_wdata_ready3;
assign hdmi2usbsoc_litedramport3_wdata_ready = controllerinjector_new_master_wdata_ready4;
assign encoder_port_port_wdata_ready = controllerinjector_new_master_wdata_ready5;
assign hdmi2usbsoc_port_rdata_valid = controllerinjector_new_master_rdata_valid5;
assign hdmi2usbsoc_litedramport0_rdata_valid0 = controllerinjector_new_master_rdata_valid11;
assign hdmi2usbsoc_litedramport1_rdata_valid0 = controllerinjector_new_master_rdata_valid17;
assign hdmi2usbsoc_litedramport2_rdata_valid0 = controllerinjector_new_master_rdata_valid23;
assign hdmi2usbsoc_litedramport3_rdata_valid0 = controllerinjector_new_master_rdata_valid29;
assign encoder_port_port_rdata_valid = controllerinjector_new_master_rdata_valid35;

// synthesis translate_off
reg dummy_d_55;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_sdram_interface_wdata <= 64'd0;
	hdmi2usbsoc_sdram_interface_wdata_we <= 8'd0;
	case ({controllerinjector_new_master_wdata_ready5, controllerinjector_new_master_wdata_ready4, controllerinjector_new_master_wdata_ready3, controllerinjector_new_master_wdata_ready2, controllerinjector_new_master_wdata_ready1, controllerinjector_new_master_wdata_ready0})
		1'd1: begin
			hdmi2usbsoc_sdram_interface_wdata <= hdmi2usbsoc_port_wdata_payload_data;
			hdmi2usbsoc_sdram_interface_wdata_we <= hdmi2usbsoc_port_wdata_payload_we;
		end
		2'd2: begin
			hdmi2usbsoc_sdram_interface_wdata <= hdmi2usbsoc_litedramport0_wdata_payload_data;
			hdmi2usbsoc_sdram_interface_wdata_we <= hdmi2usbsoc_litedramport0_wdata_payload_we;
		end
		3'd4: begin
			hdmi2usbsoc_sdram_interface_wdata <= hdmi2usbsoc_litedramport1_wdata_payload_data;
			hdmi2usbsoc_sdram_interface_wdata_we <= hdmi2usbsoc_litedramport1_wdata_payload_we;
		end
		4'd8: begin
			hdmi2usbsoc_sdram_interface_wdata <= hdmi2usbsoc_litedramport2_wdata_payload_data;
			hdmi2usbsoc_sdram_interface_wdata_we <= hdmi2usbsoc_litedramport2_wdata_payload_we;
		end
		5'd16: begin
			hdmi2usbsoc_sdram_interface_wdata <= hdmi2usbsoc_litedramport3_wdata_payload_data;
			hdmi2usbsoc_sdram_interface_wdata_we <= hdmi2usbsoc_litedramport3_wdata_payload_we;
		end
		6'd32: begin
			hdmi2usbsoc_sdram_interface_wdata <= encoder_port_port_wdata_payload_data;
			hdmi2usbsoc_sdram_interface_wdata_we <= encoder_port_port_wdata_payload_we;
		end
		default: begin
			hdmi2usbsoc_sdram_interface_wdata <= 1'd0;
			hdmi2usbsoc_sdram_interface_wdata_we <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_55 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_port_rdata_payload_data = hdmi2usbsoc_sdram_interface_rdata;
assign hdmi2usbsoc_litedramport0_rdata_payload_data0 = hdmi2usbsoc_sdram_interface_rdata;
assign hdmi2usbsoc_litedramport1_rdata_payload_data0 = hdmi2usbsoc_sdram_interface_rdata;
assign hdmi2usbsoc_litedramport2_rdata_payload_data0 = hdmi2usbsoc_sdram_interface_rdata;
assign hdmi2usbsoc_litedramport3_rdata_payload_data0 = hdmi2usbsoc_sdram_interface_rdata;
assign encoder_port_port_rdata_payload_data = hdmi2usbsoc_sdram_interface_rdata;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_din = {hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_last, hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_first, hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_payload_adr, hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_payload_we};
assign {hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_last, hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_first, hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_payload_adr, hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_payload_we} = hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_dout;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_ready = hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_writable;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_we = hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_valid;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_first = hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_first;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_last = hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_last;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_payload_we = hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_payload_we;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_in_payload_adr = hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_payload_adr;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_valid = hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_readable;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_first = hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_first;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_last = hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_last;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_payload_we = hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_payload_we;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_payload_adr = hdmi2usbsoc_litedramportcdc0_cmd_fifo_fifo_out_payload_adr;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_re = hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_ready;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_ce = (hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_writable & hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_we);
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_ce = (hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_readable & hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_re);
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_writable = (((hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q[2] == hdmi2usbsoc_litedramportcdc0_cmd_fifo_consume_wdomain[2]) | (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q[1] == hdmi2usbsoc_litedramportcdc0_cmd_fifo_consume_wdomain[1])) | (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q[0] != hdmi2usbsoc_litedramportcdc0_cmd_fifo_consume_wdomain[0]));
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_readable = (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q != hdmi2usbsoc_litedramportcdc0_cmd_fifo_produce_rdomain);
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_adr = hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_binary[1:0];
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_dat_w = hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_din;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_we = hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_ce;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_rdport_adr = hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary[1:0];
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_asyncfifo0_dout = hdmi2usbsoc_litedramportcdc0_cmd_fifo_rdport_dat_r;

// synthesis translate_off
reg dummy_d_56;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next_binary <= 3'd0;
	if (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_ce) begin
		hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next_binary <= (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next_binary <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_56 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next = (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next_binary ^ hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_57;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary <= 3'd0;
	if (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_ce) begin
		hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary <= (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_57 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next = (hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary ^ hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary[2:1]);
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_valid = hdmi2usbsoc_litedramport0_cmd_valid1;
assign hdmi2usbsoc_litedramport0_cmd_ready1 = hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_ready;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_first = hdmi2usbsoc_litedramport0_cmd_first;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_last = hdmi2usbsoc_litedramport0_cmd_last;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_payload_we = hdmi2usbsoc_litedramport0_cmd_payload_we1;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_sink_payload_adr = hdmi2usbsoc_litedramport0_cmd_payload_adr1;
assign hdmi2usbsoc_litedramport2_cmd_valid0 = hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_valid;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_ready = hdmi2usbsoc_litedramport2_cmd_ready0;
assign hdmi2usbsoc_litedramport2_cmd_first0 = hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_first;
assign hdmi2usbsoc_litedramport2_cmd_last0 = hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_last;
assign hdmi2usbsoc_litedramport2_cmd_payload_we0 = hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_payload_we;
assign hdmi2usbsoc_litedramport2_cmd_payload_adr0 = hdmi2usbsoc_litedramportcdc0_cmd_fifo_source_payload_adr;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_din = {hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_last, hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_first, hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_last, hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_first, hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_payload_data} = hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_dout;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_ready = hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_writable;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_we = hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_valid;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_first = hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_first;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_last = hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_last;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_in_payload_data = hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_payload_data;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_valid = hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_readable;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_first = hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_first;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_last = hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_last;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_payload_data = hdmi2usbsoc_litedramportcdc0_rdata_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_re = hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_ready;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_ce = (hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_writable & hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_we);
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_ce = (hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_readable & hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_re);
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_writable = (((hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q[4] == hdmi2usbsoc_litedramportcdc0_rdata_fifo_consume_wdomain[4]) | (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q[3] == hdmi2usbsoc_litedramportcdc0_rdata_fifo_consume_wdomain[3])) | (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q[2:0] != hdmi2usbsoc_litedramportcdc0_rdata_fifo_consume_wdomain[2:0]));
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_readable = (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q != hdmi2usbsoc_litedramportcdc0_rdata_fifo_produce_rdomain);
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_adr = hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_binary[3:0];
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_dat_w = hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_din;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_we = hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_ce;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_rdport_adr = hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary[3:0];
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_asyncfifo0_dout = hdmi2usbsoc_litedramportcdc0_rdata_fifo_rdport_dat_r;

// synthesis translate_off
reg dummy_d_58;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next_binary <= 5'd0;
	if (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_ce) begin
		hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next_binary <= (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next_binary <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_58 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next = (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next_binary ^ hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next_binary[4:1]);

// synthesis translate_off
reg dummy_d_59;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary <= 5'd0;
	if (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_ce) begin
		hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary <= (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_59 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next = (hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary ^ hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary[4:1]);
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_valid = hdmi2usbsoc_litedramport2_rdata_valid0;
assign hdmi2usbsoc_litedramport2_rdata_ready0 = hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_ready;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_first = hdmi2usbsoc_litedramport2_rdata_first0;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_last = hdmi2usbsoc_litedramport2_rdata_last0;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_sink_payload_data = hdmi2usbsoc_litedramport2_rdata_payload_data0;
assign hdmi2usbsoc_litedramport0_rdata_valid1 = hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_valid;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_ready = hdmi2usbsoc_litedramport0_rdata_ready;
assign hdmi2usbsoc_litedramport0_rdata_first = hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_first;
assign hdmi2usbsoc_litedramport0_rdata_last = hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_last;
assign hdmi2usbsoc_litedramport0_rdata_payload_data1 = hdmi2usbsoc_litedramportcdc0_rdata_fifo_source_payload_data;

// synthesis translate_off
reg dummy_d_60;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramport1_cmd_ready1 <= 1'd0;
	hdmi2usbsoc_litedramport0_cmd_valid1 <= 1'd0;
	hdmi2usbsoc_litedramportconverter0_counter_ce <= 1'd0;
	hdmi2usbsoc_litedramport0_cmd_payload_adr1 <= 24'd0;
	if (hdmi2usbsoc_litedramport1_cmd_valid1) begin
		if ((hdmi2usbsoc_litedramportconverter0_counter == 1'd0)) begin
			hdmi2usbsoc_litedramport0_cmd_valid1 <= 1'd1;
			hdmi2usbsoc_litedramport0_cmd_payload_adr1 <= hdmi2usbsoc_litedramport1_cmd_payload_adr1[25:2];
			hdmi2usbsoc_litedramport1_cmd_ready1 <= hdmi2usbsoc_litedramport0_cmd_ready1;
			hdmi2usbsoc_litedramportconverter0_counter_ce <= hdmi2usbsoc_litedramport0_cmd_ready1;
		end else begin
			hdmi2usbsoc_litedramport1_cmd_ready1 <= 1'd1;
			hdmi2usbsoc_litedramportconverter0_counter_ce <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_60 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_61;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_valid <= 1'd0;
	hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_payload_sel <= 4'd0;
	if ((hdmi2usbsoc_litedramport0_cmd_valid1 & hdmi2usbsoc_litedramport0_cmd_ready1)) begin
		hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_valid <= 1'd1;
		hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_payload_sel <= 4'd15;
	end
// synthesis translate_off
	dummy_d_61 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_valid = hdmi2usbsoc_litedramport0_rdata_valid1;
assign hdmi2usbsoc_litedramport0_rdata_ready = hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_ready;
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_first = hdmi2usbsoc_litedramport0_rdata_first;
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_last = hdmi2usbsoc_litedramport0_rdata_last;
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_payload_data = hdmi2usbsoc_litedramport0_rdata_payload_data1;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_valid = hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_valid;
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_ready = hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_ready;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_first = hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_first;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_last = hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_last;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_payload_data = hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_payload_data;
assign hdmi2usbsoc_litedramportconverter0_rdata_chunk_valid = ((hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_payload_sel & hdmi2usbsoc_litedramportconverter0_rdata_chunk) != 1'd0);

// synthesis translate_off
reg dummy_d_62;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramport1_rdata_valid1 <= 1'd0;
	hdmi2usbsoc_litedramport1_rdata_payload_data1 <= 16'd0;
	hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready <= 1'd0;
	if (hdmi2usbsoc_litedramport1_flush) begin
		hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready <= 1'd1;
	end else begin
		if (hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_valid) begin
			if (hdmi2usbsoc_litedramportconverter0_rdata_chunk_valid) begin
				hdmi2usbsoc_litedramport1_rdata_valid1 <= hdmi2usbsoc_litedramportconverter0_rdata_converter_source_valid;
				hdmi2usbsoc_litedramport1_rdata_payload_data1 <= hdmi2usbsoc_litedramportconverter0_rdata_converter_source_payload_data;
				hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready <= hdmi2usbsoc_litedramport1_rdata_ready;
			end else begin
				hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready <= 1'd1;
			end
		end
	end
// synthesis translate_off
	dummy_d_62 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_ready = (hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready & hdmi2usbsoc_litedramportconverter0_rdata_chunk[3]);
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_din = {hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_last, hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_first, hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_payload_sel};
assign {hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_last, hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_first, hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_payload_sel} = hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_dout;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_ready = hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_writable;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_we = hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_valid;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_first = hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_first;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_last = hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_last;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_in_payload_sel = hdmi2usbsoc_litedramportconverter0_cmd_buffer_sink_payload_sel;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_valid = hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_readable;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_first = hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_first;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_last = hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_last;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_payload_sel = hdmi2usbsoc_litedramportconverter0_cmd_buffer_fifo_out_payload_sel;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_re = hdmi2usbsoc_litedramportconverter0_cmd_buffer_source_ready;

// synthesis translate_off
reg dummy_d_63;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_litedramportconverter0_cmd_buffer_replace) begin
		hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_adr <= (hdmi2usbsoc_litedramportconverter0_cmd_buffer_produce - 1'd1);
	end else begin
		hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_adr <= hdmi2usbsoc_litedramportconverter0_cmd_buffer_produce;
	end
// synthesis translate_off
	dummy_d_63 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_dat_w = hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_din;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_we = (hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_we & (hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_writable | hdmi2usbsoc_litedramportconverter0_cmd_buffer_replace));
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_do_read = (hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_readable & hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_re);
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_rdport_adr = hdmi2usbsoc_litedramportconverter0_cmd_buffer_consume;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_dout = hdmi2usbsoc_litedramportconverter0_cmd_buffer_rdport_dat_r;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_writable = (hdmi2usbsoc_litedramportconverter0_cmd_buffer_level != 3'd4);
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_readable = (hdmi2usbsoc_litedramportconverter0_cmd_buffer_level != 1'd0);
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_pipe_ce = (hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_ready | (~hdmi2usbsoc_litedramportconverter0_rdata_buffer_valid_n));
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_ready = hdmi2usbsoc_litedramportconverter0_rdata_buffer_pipe_ce;
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_valid = hdmi2usbsoc_litedramportconverter0_rdata_buffer_valid_n;
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_busy = (1'd0 | hdmi2usbsoc_litedramportconverter0_rdata_buffer_valid_n);
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_first = hdmi2usbsoc_litedramportconverter0_rdata_buffer_first_n;
assign hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_last = hdmi2usbsoc_litedramportconverter0_rdata_buffer_last_n;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_valid = hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_valid;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_first = hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_first;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_last = hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_last;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_ready = hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_ready;

// synthesis translate_off
reg dummy_d_64;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data <= 64'd0;
	hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[15:0] <= hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_payload_data[15:0];
	hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[31:16] <= hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_payload_data[31:16];
	hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[47:32] <= hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_payload_data[47:32];
	hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[63:48] <= hdmi2usbsoc_litedramportconverter0_rdata_converter_sink_payload_data[63:48];
// synthesis translate_off
	dummy_d_64 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_valid = hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_valid;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_first = hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_first;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_last = hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_last;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_ready = hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready;
assign {hdmi2usbsoc_litedramportconverter0_rdata_converter_source_payload_data} = hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_payload_data;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_valid = hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_valid;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_ready = hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_ready;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_first = hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_first;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_last = hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_last;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_source_source_payload_data = hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_data;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_first = (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_mux == 1'd0);
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_last = (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_mux == 2'd3);
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_valid = hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_valid;
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_first = (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_first & hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_first);
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_last = (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_last & hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_last);
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_ready = (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_last & hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_ready);

// synthesis translate_off
reg dummy_d_65;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_data <= 16'd0;
	case (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_mux)
		1'd0: begin
			hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[63:48];
		end
		1'd1: begin
			hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[47:32];
		end
		2'd2: begin
			hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[31:16];
		end
		default: begin
			hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_sink_payload_data[15:0];
		end
	endcase
// synthesis translate_off
	dummy_d_65 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_payload_valid_token_count = hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_last;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_din = {hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_last, hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_first, hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_payload_adr, hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_payload_we};
assign {hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_last, hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_first, hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_payload_adr, hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_payload_we} = hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_dout;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_ready = hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_writable;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_we = hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_valid;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_first = hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_first;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_last = hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_last;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_payload_we = hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_payload_we;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_in_payload_adr = hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_payload_adr;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_valid = hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_readable;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_first = hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_first;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_last = hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_last;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_payload_we = hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_payload_we;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_payload_adr = hdmi2usbsoc_litedramportcdc1_cmd_fifo_fifo_out_payload_adr;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_re = hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_ready;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_ce = (hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_writable & hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_we);
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_ce = (hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_readable & hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_re);
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_writable = (((hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q[2] == hdmi2usbsoc_litedramportcdc1_cmd_fifo_consume_wdomain[2]) | (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q[1] == hdmi2usbsoc_litedramportcdc1_cmd_fifo_consume_wdomain[1])) | (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q[0] != hdmi2usbsoc_litedramportcdc1_cmd_fifo_consume_wdomain[0]));
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_readable = (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q != hdmi2usbsoc_litedramportcdc1_cmd_fifo_produce_rdomain);
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_adr = hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_binary[1:0];
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_dat_w = hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_din;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_we = hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_ce;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_rdport_adr = hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary[1:0];
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_asyncfifo1_dout = hdmi2usbsoc_litedramportcdc1_cmd_fifo_rdport_dat_r;

// synthesis translate_off
reg dummy_d_66;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next_binary <= 3'd0;
	if (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_ce) begin
		hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next_binary <= (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next_binary <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_66 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next = (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next_binary ^ hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_67;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary <= 3'd0;
	if (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_ce) begin
		hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary <= (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_67 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next = (hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary ^ hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary[2:1]);
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_valid = hdmi2usbsoc_litedramport2_cmd_valid1;
assign hdmi2usbsoc_litedramport2_cmd_ready1 = hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_ready;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_first = hdmi2usbsoc_litedramport2_cmd_first1;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_last = hdmi2usbsoc_litedramport2_cmd_last1;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_payload_we = hdmi2usbsoc_litedramport2_cmd_payload_we1;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_sink_payload_adr = hdmi2usbsoc_litedramport2_cmd_payload_adr1;
assign hdmi2usbsoc_litedramport3_cmd_valid0 = hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_valid;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_ready = hdmi2usbsoc_litedramport3_cmd_ready0;
assign hdmi2usbsoc_litedramport3_cmd_first = hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_first;
assign hdmi2usbsoc_litedramport3_cmd_last = hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_last;
assign hdmi2usbsoc_litedramport3_cmd_payload_we0 = hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_payload_we;
assign hdmi2usbsoc_litedramport3_cmd_payload_adr0 = hdmi2usbsoc_litedramportcdc1_cmd_fifo_source_payload_adr;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_din = {hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_last, hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_first, hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_last, hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_first, hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_payload_data} = hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_dout;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_ready = hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_writable;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_we = hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_valid;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_first = hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_first;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_last = hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_last;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_in_payload_data = hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_payload_data;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_valid = hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_readable;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_first = hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_first;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_last = hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_last;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_payload_data = hdmi2usbsoc_litedramportcdc1_rdata_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_re = hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_ready;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_ce = (hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_writable & hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_we);
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_ce = (hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_readable & hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_re);
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_writable = (((hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q[4] == hdmi2usbsoc_litedramportcdc1_rdata_fifo_consume_wdomain[4]) | (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q[3] == hdmi2usbsoc_litedramportcdc1_rdata_fifo_consume_wdomain[3])) | (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q[2:0] != hdmi2usbsoc_litedramportcdc1_rdata_fifo_consume_wdomain[2:0]));
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_readable = (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q != hdmi2usbsoc_litedramportcdc1_rdata_fifo_produce_rdomain);
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_adr = hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_binary[3:0];
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_dat_w = hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_din;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_we = hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_ce;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_rdport_adr = hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary[3:0];
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_asyncfifo1_dout = hdmi2usbsoc_litedramportcdc1_rdata_fifo_rdport_dat_r;

// synthesis translate_off
reg dummy_d_68;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next_binary <= 5'd0;
	if (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_ce) begin
		hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next_binary <= (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next_binary <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_68 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next = (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next_binary ^ hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next_binary[4:1]);

// synthesis translate_off
reg dummy_d_69;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary <= 5'd0;
	if (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_ce) begin
		hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary <= (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_69 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next = (hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary ^ hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary[4:1]);
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_valid = hdmi2usbsoc_litedramport3_rdata_valid0;
assign hdmi2usbsoc_litedramport3_rdata_ready0 = hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_ready;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_first = hdmi2usbsoc_litedramport3_rdata_first0;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_last = hdmi2usbsoc_litedramport3_rdata_last0;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_sink_payload_data = hdmi2usbsoc_litedramport3_rdata_payload_data0;
assign hdmi2usbsoc_litedramport2_rdata_valid1 = hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_valid;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_ready = hdmi2usbsoc_litedramport2_rdata_ready1;
assign hdmi2usbsoc_litedramport2_rdata_first1 = hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_first;
assign hdmi2usbsoc_litedramport2_rdata_last1 = hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_last;
assign hdmi2usbsoc_litedramport2_rdata_payload_data1 = hdmi2usbsoc_litedramportcdc1_rdata_fifo_source_payload_data;

// synthesis translate_off
reg dummy_d_70;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramport3_cmd_ready1 <= 1'd0;
	hdmi2usbsoc_litedramportconverter1_counter_ce <= 1'd0;
	hdmi2usbsoc_litedramport2_cmd_valid1 <= 1'd0;
	hdmi2usbsoc_litedramport2_cmd_payload_adr1 <= 24'd0;
	if (hdmi2usbsoc_litedramport3_cmd_valid1) begin
		if ((hdmi2usbsoc_litedramportconverter1_counter == 1'd0)) begin
			hdmi2usbsoc_litedramport2_cmd_valid1 <= 1'd1;
			hdmi2usbsoc_litedramport2_cmd_payload_adr1 <= hdmi2usbsoc_litedramport3_cmd_payload_adr1[25:2];
			hdmi2usbsoc_litedramport3_cmd_ready1 <= hdmi2usbsoc_litedramport2_cmd_ready1;
			hdmi2usbsoc_litedramportconverter1_counter_ce <= hdmi2usbsoc_litedramport2_cmd_ready1;
		end else begin
			hdmi2usbsoc_litedramport3_cmd_ready1 <= 1'd1;
			hdmi2usbsoc_litedramportconverter1_counter_ce <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_70 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_71;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_valid <= 1'd0;
	hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_payload_sel <= 4'd0;
	if ((hdmi2usbsoc_litedramport2_cmd_valid1 & hdmi2usbsoc_litedramport2_cmd_ready1)) begin
		hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_valid <= 1'd1;
		hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_payload_sel <= 4'd15;
	end
// synthesis translate_off
	dummy_d_71 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_valid = hdmi2usbsoc_litedramport2_rdata_valid1;
assign hdmi2usbsoc_litedramport2_rdata_ready1 = hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_ready;
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_first = hdmi2usbsoc_litedramport2_rdata_first1;
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_last = hdmi2usbsoc_litedramport2_rdata_last1;
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_payload_data = hdmi2usbsoc_litedramport2_rdata_payload_data1;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_valid = hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_valid;
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_ready = hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_ready;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_first = hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_first;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_last = hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_last;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_payload_data = hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_payload_data;
assign hdmi2usbsoc_litedramportconverter1_rdata_chunk_valid = ((hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_payload_sel & hdmi2usbsoc_litedramportconverter1_rdata_chunk) != 1'd0);

// synthesis translate_off
reg dummy_d_72;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready <= 1'd0;
	hdmi2usbsoc_litedramport3_rdata_payload_data1 <= 16'd0;
	hdmi2usbsoc_litedramport3_rdata_valid1 <= 1'd0;
	if (hdmi2usbsoc_litedramport3_flush) begin
		hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready <= 1'd1;
	end else begin
		if (hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_valid) begin
			if (hdmi2usbsoc_litedramportconverter1_rdata_chunk_valid) begin
				hdmi2usbsoc_litedramport3_rdata_valid1 <= hdmi2usbsoc_litedramportconverter1_rdata_converter_source_valid;
				hdmi2usbsoc_litedramport3_rdata_payload_data1 <= hdmi2usbsoc_litedramportconverter1_rdata_converter_source_payload_data;
				hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready <= hdmi2usbsoc_litedramport3_rdata_ready1;
			end else begin
				hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready <= 1'd1;
			end
		end
	end
// synthesis translate_off
	dummy_d_72 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_ready = (hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready & hdmi2usbsoc_litedramportconverter1_rdata_chunk[3]);
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_din = {hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_last, hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_first, hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_payload_sel};
assign {hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_last, hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_first, hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_payload_sel} = hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_dout;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_ready = hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_writable;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_we = hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_valid;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_first = hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_first;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_last = hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_last;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_in_payload_sel = hdmi2usbsoc_litedramportconverter1_cmd_buffer_sink_payload_sel;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_valid = hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_readable;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_first = hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_first;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_last = hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_last;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_payload_sel = hdmi2usbsoc_litedramportconverter1_cmd_buffer_fifo_out_payload_sel;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_re = hdmi2usbsoc_litedramportconverter1_cmd_buffer_source_ready;

// synthesis translate_off
reg dummy_d_73;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_litedramportconverter1_cmd_buffer_replace) begin
		hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_adr <= (hdmi2usbsoc_litedramportconverter1_cmd_buffer_produce - 1'd1);
	end else begin
		hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_adr <= hdmi2usbsoc_litedramportconverter1_cmd_buffer_produce;
	end
// synthesis translate_off
	dummy_d_73 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_dat_w = hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_din;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_we = (hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_we & (hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_writable | hdmi2usbsoc_litedramportconverter1_cmd_buffer_replace));
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_do_read = (hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_readable & hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_re);
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_rdport_adr = hdmi2usbsoc_litedramportconverter1_cmd_buffer_consume;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_dout = hdmi2usbsoc_litedramportconverter1_cmd_buffer_rdport_dat_r;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_writable = (hdmi2usbsoc_litedramportconverter1_cmd_buffer_level != 3'd4);
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_readable = (hdmi2usbsoc_litedramportconverter1_cmd_buffer_level != 1'd0);
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_pipe_ce = (hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_ready | (~hdmi2usbsoc_litedramportconverter1_rdata_buffer_valid_n));
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_ready = hdmi2usbsoc_litedramportconverter1_rdata_buffer_pipe_ce;
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_valid = hdmi2usbsoc_litedramportconverter1_rdata_buffer_valid_n;
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_busy = (1'd0 | hdmi2usbsoc_litedramportconverter1_rdata_buffer_valid_n);
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_first = hdmi2usbsoc_litedramportconverter1_rdata_buffer_first_n;
assign hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_last = hdmi2usbsoc_litedramportconverter1_rdata_buffer_last_n;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_valid = hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_valid;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_first = hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_first;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_last = hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_last;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_ready = hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_ready;

// synthesis translate_off
reg dummy_d_74;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data <= 64'd0;
	hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[15:0] <= hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_payload_data[15:0];
	hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[31:16] <= hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_payload_data[31:16];
	hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[47:32] <= hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_payload_data[47:32];
	hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[63:48] <= hdmi2usbsoc_litedramportconverter1_rdata_converter_sink_payload_data[63:48];
// synthesis translate_off
	dummy_d_74 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_valid = hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_valid;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_first = hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_first;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_last = hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_last;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_ready = hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready;
assign {hdmi2usbsoc_litedramportconverter1_rdata_converter_source_payload_data} = hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_payload_data;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_valid = hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_valid;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_ready = hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_ready;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_first = hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_first;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_last = hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_last;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_source_source_payload_data = hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_data;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_first = (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_mux == 1'd0);
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_last = (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_mux == 2'd3);
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_valid = hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_valid;
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_first = (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_first & hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_first);
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_last = (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_last & hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_last);
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_ready = (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_last & hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_ready);

// synthesis translate_off
reg dummy_d_75;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_data <= 16'd0;
	case (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_mux)
		1'd0: begin
			hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[63:48];
		end
		1'd1: begin
			hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[47:32];
		end
		2'd2: begin
			hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[31:16];
		end
		default: begin
			hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_data <= hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_sink_payload_data[15:0];
		end
	endcase
// synthesis translate_off
	dummy_d_75 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_payload_valid_token_count = hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_last;

// synthesis translate_off
reg dummy_d_76;
// synthesis translate_on
always @(*) begin
	controllerinjector_next_state <= 1'd0;
	encoder_port_port_cmd_valid <= 1'd0;
	encoder_port_port_cmd_payload_we <= 1'd0;
	encoder_port_new_port_cmd_ready <= 1'd0;
	encoder_port_port_cmd_payload_adr <= 24'd0;
	encoder_port_counter_reset <= 1'd0;
	encoder_port_counter_ce <= 1'd0;
	controllerinjector_next_state <= controllerinjector_state;
	case (controllerinjector_state)
		1'd1: begin
			encoder_port_port_cmd_valid <= 1'd1;
			encoder_port_port_cmd_payload_we <= encoder_port_new_port_cmd_payload_we;
			encoder_port_port_cmd_payload_adr <= ((encoder_port_new_port_cmd_payload_adr * 2'd2) + encoder_port_counter);
			if (encoder_port_port_cmd_ready) begin
				encoder_port_counter_ce <= 1'd1;
				if ((encoder_port_counter == 1'd1)) begin
					encoder_port_new_port_cmd_ready <= 1'd1;
					controllerinjector_next_state <= 1'd0;
				end
			end
		end
		default: begin
			encoder_port_counter_reset <= 1'd1;
			if (encoder_port_new_port_cmd_valid) begin
				controllerinjector_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_76 <= dummy_s;
// synthesis translate_on
end
assign encoder_port_converter_sink_valid = encoder_port_sink_valid;
assign encoder_port_converter_sink_first = encoder_port_sink_first;
assign encoder_port_converter_sink_last = encoder_port_sink_last;
assign encoder_port_sink_ready = encoder_port_converter_sink_ready;
assign encoder_port_converter_sink_payload_data = {encoder_port_sink_payload_data};
assign encoder_port_source_valid = encoder_port_source_source_valid;
assign encoder_port_source_first = encoder_port_source_source_first;
assign encoder_port_source_last = encoder_port_source_source_last;
assign encoder_port_source_source_ready = encoder_port_source_ready;

// synthesis translate_off
reg dummy_d_77;
// synthesis translate_on
always @(*) begin
	encoder_port_source_payload_data <= 128'd0;
	encoder_port_source_payload_data[63:0] <= encoder_port_source_source_payload_data[63:0];
	encoder_port_source_payload_data[127:64] <= encoder_port_source_source_payload_data[127:64];
// synthesis translate_off
	dummy_d_77 <= dummy_s;
// synthesis translate_on
end
assign encoder_port_source_source_valid = encoder_port_converter_source_valid;
assign encoder_port_converter_source_ready = encoder_port_source_source_ready;
assign encoder_port_source_source_first = encoder_port_converter_source_first;
assign encoder_port_source_source_last = encoder_port_converter_source_last;
assign encoder_port_source_source_payload_data = encoder_port_converter_source_payload_data;
assign encoder_port_converter_sink_ready = ((~encoder_port_converter_strobe_all) | encoder_port_converter_source_ready);
assign encoder_port_converter_source_valid = encoder_port_converter_strobe_all;
assign encoder_port_converter_load_part = (encoder_port_converter_sink_valid & encoder_port_converter_sink_ready);
assign encoder_port_sink_valid = encoder_port_port_rdata_valid;
assign encoder_port_port_rdata_ready = encoder_port_sink_ready;
assign encoder_port_sink_first = encoder_port_port_rdata_first;
assign encoder_port_sink_last = encoder_port_port_rdata_last;
assign encoder_port_sink_payload_data = encoder_port_port_rdata_payload_data;
assign encoder_port_new_port_rdata_valid = encoder_port_source_valid;
assign encoder_port_source_ready = encoder_port_new_port_rdata_ready;
assign encoder_port_new_port_rdata_first = encoder_port_source_first;
assign encoder_port_new_port_rdata_last = encoder_port_source_last;
assign encoder_port_new_port_rdata_payload_data = encoder_port_source_payload_data;
assign hdmi2usbsoc_data_port_adr = hdmi2usbsoc_interface0_wb_sdram_adr[10:1];

// synthesis translate_off
reg dummy_d_78;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_data_port_dat_w <= 64'd0;
	hdmi2usbsoc_data_port_we <= 8'd0;
	if (hdmi2usbsoc_write_from_slave) begin
		hdmi2usbsoc_data_port_dat_w <= hdmi2usbsoc_interface_dat_r;
		hdmi2usbsoc_data_port_we <= {8{1'd1}};
	end else begin
		hdmi2usbsoc_data_port_dat_w <= {2{hdmi2usbsoc_interface0_wb_sdram_dat_w}};
		if ((((hdmi2usbsoc_interface0_wb_sdram_cyc & hdmi2usbsoc_interface0_wb_sdram_stb) & hdmi2usbsoc_interface0_wb_sdram_we) & hdmi2usbsoc_interface0_wb_sdram_ack)) begin
			hdmi2usbsoc_data_port_we <= {({4{(hdmi2usbsoc_interface0_wb_sdram_adr[0] == 1'd0)}} & hdmi2usbsoc_interface0_wb_sdram_sel), ({4{(hdmi2usbsoc_interface0_wb_sdram_adr[0] == 1'd1)}} & hdmi2usbsoc_interface0_wb_sdram_sel)};
		end
	end
// synthesis translate_off
	dummy_d_78 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_interface_dat_w = hdmi2usbsoc_data_port_dat_r;
assign hdmi2usbsoc_interface_sel = 8'd255;

// synthesis translate_off
reg dummy_d_79;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_interface0_wb_sdram_dat_r <= 32'd0;
	case (hdmi2usbsoc_adr_offset_r)
		1'd0: begin
			hdmi2usbsoc_interface0_wb_sdram_dat_r <= hdmi2usbsoc_data_port_dat_r[63:32];
		end
		default: begin
			hdmi2usbsoc_interface0_wb_sdram_dat_r <= hdmi2usbsoc_data_port_dat_r[31:0];
		end
	endcase
// synthesis translate_off
	dummy_d_79 <= dummy_s;
// synthesis translate_on
end
assign {hdmi2usbsoc_tag_do_dirty, hdmi2usbsoc_tag_do_tag} = hdmi2usbsoc_tag_port_dat_r;
assign hdmi2usbsoc_tag_port_dat_w = {hdmi2usbsoc_tag_di_dirty, hdmi2usbsoc_tag_di_tag};
assign hdmi2usbsoc_tag_port_adr = hdmi2usbsoc_interface0_wb_sdram_adr[10:1];
assign hdmi2usbsoc_tag_di_tag = hdmi2usbsoc_interface0_wb_sdram_adr[29:11];
assign hdmi2usbsoc_interface_adr = {hdmi2usbsoc_tag_do_tag, hdmi2usbsoc_interface0_wb_sdram_adr[10:1]};

// synthesis translate_off
reg dummy_d_80;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_tag_port_we <= 1'd0;
	hdmi2usbsoc_interface_cyc <= 1'd0;
	hdmi2usbsoc_interface_stb <= 1'd0;
	hdmi2usbsoc_tag_di_dirty <= 1'd0;
	hdmi2usbsoc_interface_we <= 1'd0;
	hdmi2usbsoc_word_clr <= 1'd0;
	hdmi2usbsoc_word_inc <= 1'd0;
	cache_next_state <= 3'd0;
	hdmi2usbsoc_interface0_wb_sdram_ack <= 1'd0;
	hdmi2usbsoc_write_from_slave <= 1'd0;
	cache_next_state <= cache_state;
	case (cache_state)
		1'd1: begin
			hdmi2usbsoc_word_clr <= 1'd1;
			if ((hdmi2usbsoc_tag_do_tag == hdmi2usbsoc_interface0_wb_sdram_adr[29:11])) begin
				hdmi2usbsoc_interface0_wb_sdram_ack <= 1'd1;
				if (hdmi2usbsoc_interface0_wb_sdram_we) begin
					hdmi2usbsoc_tag_di_dirty <= 1'd1;
					hdmi2usbsoc_tag_port_we <= 1'd1;
				end
				cache_next_state <= 1'd0;
			end else begin
				if (hdmi2usbsoc_tag_do_dirty) begin
					cache_next_state <= 2'd2;
				end else begin
					cache_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			hdmi2usbsoc_interface_stb <= 1'd1;
			hdmi2usbsoc_interface_cyc <= 1'd1;
			hdmi2usbsoc_interface_we <= 1'd1;
			if (hdmi2usbsoc_interface_ack) begin
				hdmi2usbsoc_word_inc <= 1'd1;
				if (1'd1) begin
					cache_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			hdmi2usbsoc_tag_port_we <= 1'd1;
			hdmi2usbsoc_word_clr <= 1'd1;
			cache_next_state <= 3'd4;
		end
		3'd4: begin
			hdmi2usbsoc_interface_stb <= 1'd1;
			hdmi2usbsoc_interface_cyc <= 1'd1;
			hdmi2usbsoc_interface_we <= 1'd0;
			if (hdmi2usbsoc_interface_ack) begin
				hdmi2usbsoc_write_from_slave <= 1'd1;
				hdmi2usbsoc_word_inc <= 1'd1;
				if (1'd1) begin
					cache_next_state <= 1'd1;
				end else begin
					cache_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((hdmi2usbsoc_interface0_wb_sdram_cyc & hdmi2usbsoc_interface0_wb_sdram_stb)) begin
				cache_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_80 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_port_cmd_payload_adr = hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_port_wdata_payload_we = hdmi2usbsoc_interface_sel;
assign hdmi2usbsoc_port_wdata_payload_data = hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface_dat_r = hdmi2usbsoc_port_rdata_payload_data;

// synthesis translate_off
reg dummy_d_81;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_port_rdata_ready <= 1'd0;
	hdmi2usbsoc_port_cmd_valid <= 1'd0;
	hdmi2usbsoc_port_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_port_wdata_valid <= 1'd0;
	hdmi2usbsoc_interface_ack <= 1'd0;
	litedramwishbonebridge_next_state <= 2'd0;
	litedramwishbonebridge_next_state <= litedramwishbonebridge_state;
	case (litedramwishbonebridge_state)
		1'd1: begin
			hdmi2usbsoc_port_cmd_valid <= 1'd1;
			hdmi2usbsoc_port_cmd_payload_we <= hdmi2usbsoc_interface_we;
			if (hdmi2usbsoc_port_cmd_ready) begin
				if (hdmi2usbsoc_interface_we) begin
					litedramwishbonebridge_next_state <= 2'd2;
				end else begin
					litedramwishbonebridge_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			hdmi2usbsoc_port_wdata_valid <= 1'd1;
			if (hdmi2usbsoc_port_wdata_ready) begin
				hdmi2usbsoc_interface_ack <= 1'd1;
				litedramwishbonebridge_next_state <= 1'd0;
			end
		end
		2'd3: begin
			hdmi2usbsoc_port_rdata_ready <= 1'd1;
			if (hdmi2usbsoc_port_rdata_valid) begin
				hdmi2usbsoc_interface_ack <= 1'd1;
				litedramwishbonebridge_next_state <= 1'd0;
			end
		end
		default: begin
			if ((hdmi2usbsoc_interface_cyc & hdmi2usbsoc_interface_stb)) begin
				litedramwishbonebridge_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_81 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_serdesstrobe = hdmi2usbsoc_hdmi_in0_serdesstrobe;
assign hdmi2usbsoc_hdmi_in0_charsync0_raw_data = hdmi2usbsoc_hdmi_in0_s6datacapture0_d;
assign hdmi2usbsoc_hdmi_in0_wer0_data = hdmi2usbsoc_hdmi_in0_charsync0_data;
assign hdmi2usbsoc_hdmi_in0_decoding0_valid_i = hdmi2usbsoc_hdmi_in0_charsync0_synced;
assign hdmi2usbsoc_hdmi_in0_decoding0_input = hdmi2usbsoc_hdmi_in0_charsync0_data;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_serdesstrobe = hdmi2usbsoc_hdmi_in0_serdesstrobe;
assign hdmi2usbsoc_hdmi_in0_charsync1_raw_data = hdmi2usbsoc_hdmi_in0_s6datacapture1_d;
assign hdmi2usbsoc_hdmi_in0_wer1_data = hdmi2usbsoc_hdmi_in0_charsync1_data;
assign hdmi2usbsoc_hdmi_in0_decoding1_valid_i = hdmi2usbsoc_hdmi_in0_charsync1_synced;
assign hdmi2usbsoc_hdmi_in0_decoding1_input = hdmi2usbsoc_hdmi_in0_charsync1_data;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_serdesstrobe = hdmi2usbsoc_hdmi_in0_serdesstrobe;
assign hdmi2usbsoc_hdmi_in0_charsync2_raw_data = hdmi2usbsoc_hdmi_in0_s6datacapture2_d;
assign hdmi2usbsoc_hdmi_in0_wer2_data = hdmi2usbsoc_hdmi_in0_charsync2_data;
assign hdmi2usbsoc_hdmi_in0_decoding2_valid_i = hdmi2usbsoc_hdmi_in0_charsync2_synced;
assign hdmi2usbsoc_hdmi_in0_decoding2_input = hdmi2usbsoc_hdmi_in0_charsync2_data;
assign hdmi2usbsoc_hdmi_in0_chansync_valid_i = ((hdmi2usbsoc_hdmi_in0_decoding0_valid_o & hdmi2usbsoc_hdmi_in0_decoding1_valid_o) & hdmi2usbsoc_hdmi_in0_decoding2_valid_o);
assign hdmi2usbsoc_hdmi_in0_chansync_data_in0_raw = hdmi2usbsoc_hdmi_in0_decoding0_output_raw;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in0_d = hdmi2usbsoc_hdmi_in0_decoding0_output_d;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in0_c = hdmi2usbsoc_hdmi_in0_decoding0_output_c;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in0_de = hdmi2usbsoc_hdmi_in0_decoding0_output_de;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in1_raw = hdmi2usbsoc_hdmi_in0_decoding1_output_raw;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in1_d = hdmi2usbsoc_hdmi_in0_decoding1_output_d;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in1_c = hdmi2usbsoc_hdmi_in0_decoding1_output_c;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in1_de = hdmi2usbsoc_hdmi_in0_decoding1_output_de;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in2_raw = hdmi2usbsoc_hdmi_in0_decoding2_output_raw;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in2_d = hdmi2usbsoc_hdmi_in0_decoding2_output_d;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in2_c = hdmi2usbsoc_hdmi_in0_decoding2_output_c;
assign hdmi2usbsoc_hdmi_in0_chansync_data_in2_de = hdmi2usbsoc_hdmi_in0_decoding2_output_de;
assign hdmi2usbsoc_hdmi_in0_syncpol_valid_i = hdmi2usbsoc_hdmi_in0_chansync_chan_synced;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in0_raw = hdmi2usbsoc_hdmi_in0_chansync_data_out0_raw;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in0_d = hdmi2usbsoc_hdmi_in0_chansync_data_out0_d;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in0_c = hdmi2usbsoc_hdmi_in0_chansync_data_out0_c;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in0_de = hdmi2usbsoc_hdmi_in0_chansync_data_out0_de;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in1_raw = hdmi2usbsoc_hdmi_in0_chansync_data_out1_raw;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in1_d = hdmi2usbsoc_hdmi_in0_chansync_data_out1_d;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in1_c = hdmi2usbsoc_hdmi_in0_chansync_data_out1_c;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in1_de = hdmi2usbsoc_hdmi_in0_chansync_data_out1_de;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in2_raw = hdmi2usbsoc_hdmi_in0_chansync_data_out2_raw;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in2_d = hdmi2usbsoc_hdmi_in0_chansync_data_out2_d;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in2_c = hdmi2usbsoc_hdmi_in0_chansync_data_out2_c;
assign hdmi2usbsoc_hdmi_in0_syncpol_data_in2_de = hdmi2usbsoc_hdmi_in0_chansync_data_out2_de;
assign hdmi2usbsoc_hdmi_in0_resdetection_valid_i = hdmi2usbsoc_hdmi_in0_syncpol_valid_o;
assign hdmi2usbsoc_hdmi_in0_resdetection_de = hdmi2usbsoc_hdmi_in0_syncpol_de;
assign hdmi2usbsoc_hdmi_in0_resdetection_vsync = hdmi2usbsoc_hdmi_in0_syncpol_vsync;
assign hdmi2usbsoc_hdmi_in0_frame_valid_i = hdmi2usbsoc_hdmi_in0_syncpol_valid_o;
assign hdmi2usbsoc_hdmi_in0_frame_de = hdmi2usbsoc_hdmi_in0_syncpol_de;
assign hdmi2usbsoc_hdmi_in0_frame_vsync = hdmi2usbsoc_hdmi_in0_syncpol_vsync;
assign hdmi2usbsoc_hdmi_in0_frame_r = hdmi2usbsoc_hdmi_in0_syncpol_r;
assign hdmi2usbsoc_hdmi_in0_frame_g = hdmi2usbsoc_hdmi_in0_syncpol_g;
assign hdmi2usbsoc_hdmi_in0_frame_b = hdmi2usbsoc_hdmi_in0_syncpol_b;
assign hdmi2usbsoc_hdmi_in0_dma_frame_valid = hdmi2usbsoc_hdmi_in0_frame_frame_valid;
assign hdmi2usbsoc_hdmi_in0_frame_frame_ready = hdmi2usbsoc_hdmi_in0_dma_frame_ready;
assign hdmi2usbsoc_hdmi_in0_dma_frame_first = hdmi2usbsoc_hdmi_in0_frame_frame_first;
assign hdmi2usbsoc_hdmi_in0_dma_frame_last = hdmi2usbsoc_hdmi_in0_frame_frame_last;
assign hdmi2usbsoc_hdmi_in0_dma_frame_payload_sof = hdmi2usbsoc_hdmi_in0_frame_frame_payload_sof;
assign hdmi2usbsoc_hdmi_in0_dma_frame_payload_pixels = hdmi2usbsoc_hdmi_in0_frame_frame_payload_pixels;
assign hdmi2usbsoc_hdmi_in0_edid_status = 1'd1;
assign hdmi2usbsoc_hdmi_in0_edid_sda_o = (~hdmi2usbsoc_hdmi_in0_edid_sda_drv_reg);
assign hdmi2usbsoc_hdmi_in0_edid_scl_rising = (hdmi2usbsoc_hdmi_in0_edid_scl_i & (~hdmi2usbsoc_hdmi_in0_edid_scl_r));
assign hdmi2usbsoc_hdmi_in0_edid_sda_rising = (hdmi2usbsoc_hdmi_in0_edid_sda_i & (~hdmi2usbsoc_hdmi_in0_edid_sda_r));
assign hdmi2usbsoc_hdmi_in0_edid_sda_falling = ((~hdmi2usbsoc_hdmi_in0_edid_sda_i) & hdmi2usbsoc_hdmi_in0_edid_sda_r);
assign hdmi2usbsoc_hdmi_in0_edid_start = (hdmi2usbsoc_hdmi_in0_edid_scl_i & hdmi2usbsoc_hdmi_in0_edid_sda_falling);
assign hdmi2usbsoc_hdmi_in0_edid_adr = hdmi2usbsoc_hdmi_in0_edid_offset_counter;

// synthesis translate_off
reg dummy_d_82;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_edid_sda_drv <= 1'd0;
	if (hdmi2usbsoc_hdmi_in0_edid_zero_drv) begin
		hdmi2usbsoc_hdmi_in0_edid_sda_drv <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_edid_data_drv) begin
			hdmi2usbsoc_hdmi_in0_edid_sda_drv <= (~hdmi2usbsoc_hdmi_in0_edid_data_bit);
		end
	end
// synthesis translate_off
	dummy_d_82 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_83;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_edid_update_is_read <= 1'd0;
	hdmi2usbsoc_hdmi_in0_edid_oc_load <= 1'd0;
	hdmi2usbsoc_hdmi_in0_edid_oc_inc <= 1'd0;
	edid0_next_state <= 4'd0;
	hdmi2usbsoc_hdmi_in0_edid_zero_drv <= 1'd0;
	hdmi2usbsoc_hdmi_in0_edid_data_drv_en <= 1'd0;
	hdmi2usbsoc_hdmi_in0_edid_data_drv_stop <= 1'd0;
	edid0_next_state <= edid0_state;
	case (edid0_state)
		1'd1: begin
			if ((hdmi2usbsoc_hdmi_in0_edid_counter == 4'd8)) begin
				if ((hdmi2usbsoc_hdmi_in0_edid_din[7:1] == 7'd80)) begin
					hdmi2usbsoc_hdmi_in0_edid_update_is_read <= 1'd1;
					edid0_next_state <= 2'd2;
				end else begin
					edid0_next_state <= 1'd0;
				end
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		2'd2: begin
			if ((~hdmi2usbsoc_hdmi_in0_edid_scl_i)) begin
				edid0_next_state <= 2'd3;
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		2'd3: begin
			hdmi2usbsoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if (hdmi2usbsoc_hdmi_in0_edid_scl_i) begin
				edid0_next_state <= 3'd4;
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		3'd4: begin
			hdmi2usbsoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if ((~hdmi2usbsoc_hdmi_in0_edid_scl_i)) begin
				if (hdmi2usbsoc_hdmi_in0_edid_is_read) begin
					edid0_next_state <= 4'd9;
				end else begin
					edid0_next_state <= 3'd5;
				end
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		3'd5: begin
			if ((hdmi2usbsoc_hdmi_in0_edid_counter == 4'd8)) begin
				hdmi2usbsoc_hdmi_in0_edid_oc_load <= 1'd1;
				edid0_next_state <= 3'd6;
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		3'd6: begin
			if ((~hdmi2usbsoc_hdmi_in0_edid_scl_i)) begin
				edid0_next_state <= 3'd7;
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		3'd7: begin
			hdmi2usbsoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if (hdmi2usbsoc_hdmi_in0_edid_scl_i) begin
				edid0_next_state <= 4'd8;
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		4'd8: begin
			hdmi2usbsoc_hdmi_in0_edid_zero_drv <= 1'd1;
			if ((~hdmi2usbsoc_hdmi_in0_edid_scl_i)) begin
				edid0_next_state <= 1'd1;
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		4'd9: begin
			if ((~hdmi2usbsoc_hdmi_in0_edid_scl_i)) begin
				if ((hdmi2usbsoc_hdmi_in0_edid_counter == 4'd8)) begin
					hdmi2usbsoc_hdmi_in0_edid_data_drv_stop <= 1'd1;
					edid0_next_state <= 4'd10;
				end else begin
					hdmi2usbsoc_hdmi_in0_edid_data_drv_en <= 1'd1;
				end
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		4'd10: begin
			if (hdmi2usbsoc_hdmi_in0_edid_scl_rising) begin
				hdmi2usbsoc_hdmi_in0_edid_oc_inc <= 1'd1;
				if (hdmi2usbsoc_hdmi_in0_edid_sda_i) begin
					edid0_next_state <= 1'd0;
				end else begin
					edid0_next_state <= 4'd9;
				end
			end
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
		default: begin
			if (hdmi2usbsoc_hdmi_in0_edid_start) begin
				edid0_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_83 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_locked_status = hdmi2usbsoc_hdmi_in0_locked;
assign hdmi_in0_pix_o_clk = hdmi_in0_pix_clk;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_too_late = (hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness == 8'd255);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_too_early = (hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness == 1'd0);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_cal = hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_rst = hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_cal = hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_rst = hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_inc = hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_ce = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_o | hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_o);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_i = (hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r[0]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_i = (hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r[1]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_i = (hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r[2]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_i = (hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r[3]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_i = (hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r[4]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_i = (hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r[5]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_busy_status = {hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_slave_pending, hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_master_pending};
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_reset_lateness = hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_i = hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_reset_re;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_o = (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_charsync0_raw = {hdmi2usbsoc_hdmi_in0_charsync0_raw_data, hdmi2usbsoc_hdmi_in0_charsync0_raw_data1};

// synthesis translate_off
reg dummy_d_84;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_wer0_transitions <= 8'd0;
	hdmi2usbsoc_hdmi_in0_wer0_transitions[0] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[0] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[1]);
	hdmi2usbsoc_hdmi_in0_wer0_transitions[1] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[1] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[2]);
	hdmi2usbsoc_hdmi_in0_wer0_transitions[2] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[2] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[3]);
	hdmi2usbsoc_hdmi_in0_wer0_transitions[3] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[3] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[4]);
	hdmi2usbsoc_hdmi_in0_wer0_transitions[4] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[4] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[5]);
	hdmi2usbsoc_hdmi_in0_wer0_transitions[5] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[5] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[6]);
	hdmi2usbsoc_hdmi_in0_wer0_transitions[6] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[6] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[7]);
	hdmi2usbsoc_hdmi_in0_wer0_transitions[7] <= (hdmi2usbsoc_hdmi_in0_wer0_data_r[7] ^ hdmi2usbsoc_hdmi_in0_wer0_data_r[8]);
// synthesis translate_off
	dummy_d_84 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_wer0_i = hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r_updated;
assign hdmi2usbsoc_hdmi_in0_wer0_o = (hdmi2usbsoc_hdmi_in0_wer0_toggle_o ^ hdmi2usbsoc_hdmi_in0_wer0_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_too_late = (hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness == 8'd255);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_too_early = (hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness == 1'd0);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_cal = hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_rst = hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_cal = hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_rst = hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_inc = hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_ce = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_o | hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_o);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_i = (hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r[0]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_i = (hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r[1]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_i = (hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r[2]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_i = (hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r[3]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_i = (hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r[4]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_i = (hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r[5]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_busy_status = {hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_slave_pending, hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_master_pending};
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_reset_lateness = hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_i = hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_reset_re;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_o = (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_charsync1_raw = {hdmi2usbsoc_hdmi_in0_charsync1_raw_data, hdmi2usbsoc_hdmi_in0_charsync1_raw_data1};

// synthesis translate_off
reg dummy_d_85;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_wer1_transitions <= 8'd0;
	hdmi2usbsoc_hdmi_in0_wer1_transitions[0] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[0] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[1]);
	hdmi2usbsoc_hdmi_in0_wer1_transitions[1] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[1] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[2]);
	hdmi2usbsoc_hdmi_in0_wer1_transitions[2] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[2] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[3]);
	hdmi2usbsoc_hdmi_in0_wer1_transitions[3] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[3] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[4]);
	hdmi2usbsoc_hdmi_in0_wer1_transitions[4] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[4] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[5]);
	hdmi2usbsoc_hdmi_in0_wer1_transitions[5] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[5] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[6]);
	hdmi2usbsoc_hdmi_in0_wer1_transitions[6] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[6] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[7]);
	hdmi2usbsoc_hdmi_in0_wer1_transitions[7] <= (hdmi2usbsoc_hdmi_in0_wer1_data_r[7] ^ hdmi2usbsoc_hdmi_in0_wer1_data_r[8]);
// synthesis translate_off
	dummy_d_85 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_wer1_i = hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r_updated;
assign hdmi2usbsoc_hdmi_in0_wer1_o = (hdmi2usbsoc_hdmi_in0_wer1_toggle_o ^ hdmi2usbsoc_hdmi_in0_wer1_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_too_late = (hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness == 8'd255);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_too_early = (hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness == 1'd0);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_cal = hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_rst = hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_cal = hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_rst = hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_inc = hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_ce = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_o | hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_o);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_i = (hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r[0]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_i = (hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r[1]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_i = (hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r[2]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_i = (hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r[3]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_i = (hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r[4]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_i = (hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r[5]);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_busy_status = {hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_slave_pending, hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_master_pending};
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_reset_lateness = hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_o;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_i = hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_reset_re;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_o = (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_o ^ hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_charsync2_raw = {hdmi2usbsoc_hdmi_in0_charsync2_raw_data, hdmi2usbsoc_hdmi_in0_charsync2_raw_data1};

// synthesis translate_off
reg dummy_d_86;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_wer2_transitions <= 8'd0;
	hdmi2usbsoc_hdmi_in0_wer2_transitions[0] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[0] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[1]);
	hdmi2usbsoc_hdmi_in0_wer2_transitions[1] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[1] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[2]);
	hdmi2usbsoc_hdmi_in0_wer2_transitions[2] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[2] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[3]);
	hdmi2usbsoc_hdmi_in0_wer2_transitions[3] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[3] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[4]);
	hdmi2usbsoc_hdmi_in0_wer2_transitions[4] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[4] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[5]);
	hdmi2usbsoc_hdmi_in0_wer2_transitions[5] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[5] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[6]);
	hdmi2usbsoc_hdmi_in0_wer2_transitions[6] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[6] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[7]);
	hdmi2usbsoc_hdmi_in0_wer2_transitions[7] <= (hdmi2usbsoc_hdmi_in0_wer2_data_r[7] ^ hdmi2usbsoc_hdmi_in0_wer2_data_r[8]);
// synthesis translate_off
	dummy_d_86 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_wer2_i = hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r_updated;
assign hdmi2usbsoc_hdmi_in0_wer2_o = (hdmi2usbsoc_hdmi_in0_wer2_toggle_o ^ hdmi2usbsoc_hdmi_in0_wer2_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_din = {hdmi2usbsoc_hdmi_in0_chansync_data_in0_de, hdmi2usbsoc_hdmi_in0_chansync_data_in0_c, hdmi2usbsoc_hdmi_in0_chansync_data_in0_d, hdmi2usbsoc_hdmi_in0_chansync_data_in0_raw};
assign {hdmi2usbsoc_hdmi_in0_chansync_data_out0_de, hdmi2usbsoc_hdmi_in0_chansync_data_out0_c, hdmi2usbsoc_hdmi_in0_chansync_data_out0_d, hdmi2usbsoc_hdmi_in0_chansync_data_out0_raw} = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_dout;
assign hdmi2usbsoc_hdmi_in0_chansync_is_control0 = (~hdmi2usbsoc_hdmi_in0_chansync_data_out0_de);
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_re = ((~hdmi2usbsoc_hdmi_in0_chansync_is_control0) | hdmi2usbsoc_hdmi_in0_chansync_all_control);
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_din = {hdmi2usbsoc_hdmi_in0_chansync_data_in1_de, hdmi2usbsoc_hdmi_in0_chansync_data_in1_c, hdmi2usbsoc_hdmi_in0_chansync_data_in1_d, hdmi2usbsoc_hdmi_in0_chansync_data_in1_raw};
assign {hdmi2usbsoc_hdmi_in0_chansync_data_out1_de, hdmi2usbsoc_hdmi_in0_chansync_data_out1_c, hdmi2usbsoc_hdmi_in0_chansync_data_out1_d, hdmi2usbsoc_hdmi_in0_chansync_data_out1_raw} = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_dout;
assign hdmi2usbsoc_hdmi_in0_chansync_is_control1 = (~hdmi2usbsoc_hdmi_in0_chansync_data_out1_de);
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_re = ((~hdmi2usbsoc_hdmi_in0_chansync_is_control1) | hdmi2usbsoc_hdmi_in0_chansync_all_control);
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_din = {hdmi2usbsoc_hdmi_in0_chansync_data_in2_de, hdmi2usbsoc_hdmi_in0_chansync_data_in2_c, hdmi2usbsoc_hdmi_in0_chansync_data_in2_d, hdmi2usbsoc_hdmi_in0_chansync_data_in2_raw};
assign {hdmi2usbsoc_hdmi_in0_chansync_data_out2_de, hdmi2usbsoc_hdmi_in0_chansync_data_out2_c, hdmi2usbsoc_hdmi_in0_chansync_data_out2_d, hdmi2usbsoc_hdmi_in0_chansync_data_out2_raw} = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_dout;
assign hdmi2usbsoc_hdmi_in0_chansync_is_control2 = (~hdmi2usbsoc_hdmi_in0_chansync_data_out2_de);
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_re = ((~hdmi2usbsoc_hdmi_in0_chansync_is_control2) | hdmi2usbsoc_hdmi_in0_chansync_all_control);
assign hdmi2usbsoc_hdmi_in0_chansync_all_control = ((hdmi2usbsoc_hdmi_in0_chansync_is_control0 & hdmi2usbsoc_hdmi_in0_chansync_is_control1) & hdmi2usbsoc_hdmi_in0_chansync_is_control2);
assign hdmi2usbsoc_hdmi_in0_chansync_some_control = ((hdmi2usbsoc_hdmi_in0_chansync_is_control0 | hdmi2usbsoc_hdmi_in0_chansync_is_control1) | hdmi2usbsoc_hdmi_in0_chansync_is_control2);
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_adr = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_produce;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_w = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_din;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_we = 1'd1;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_rdport_adr = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_consume;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_dout = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_adr = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_produce;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_w = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_din;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_we = 1'd1;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_rdport_adr = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_consume;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_dout = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_adr = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_produce;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_w = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_din;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_we = 1'd1;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_rdport_adr = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_consume;
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_dout = hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in0_syncpol_de = hdmi2usbsoc_hdmi_in0_syncpol_de_r;
assign hdmi2usbsoc_hdmi_in0_syncpol_hsync = hdmi2usbsoc_hdmi_in0_syncpol_c_out[0];
assign hdmi2usbsoc_hdmi_in0_syncpol_vsync = hdmi2usbsoc_hdmi_in0_syncpol_c_out[1];
assign hdmi2usbsoc_hdmi_in0_resdetection_pn_de = ((~hdmi2usbsoc_hdmi_in0_resdetection_de) & hdmi2usbsoc_hdmi_in0_resdetection_de_r);
assign hdmi2usbsoc_hdmi_in0_resdetection_p_vsync = (hdmi2usbsoc_hdmi_in0_resdetection_vsync & (~hdmi2usbsoc_hdmi_in0_resdetection_vsync_r));
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_valid = hdmi2usbsoc_hdmi_in0_frame_valid_i;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_r = hdmi2usbsoc_hdmi_in0_frame_r;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_g = hdmi2usbsoc_hdmi_in0_frame_g;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_b = hdmi2usbsoc_hdmi_in0_frame_b;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_valid = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_valid;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_ready = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_ready;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_first = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_first;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_last = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_last;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_y = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_y;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_cb = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_cb;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_cr = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_cr;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_ready = 1'd1;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first = (hdmi2usbsoc_hdmi_in0_frame_de & (~hdmi2usbsoc_hdmi_in0_frame_de_r));
assign hdmi2usbsoc_hdmi_in0_frame_new_frame = (hdmi2usbsoc_hdmi_in0_frame_next_vsync10 & (~hdmi2usbsoc_hdmi_in0_frame_vsync_r));
assign hdmi2usbsoc_hdmi_in0_frame_encoded_pixel = {hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_payload_cb_cr, hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_payload_y};
assign hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_pixels = hdmi2usbsoc_hdmi_in0_frame_cur_word;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_sink_valid = hdmi2usbsoc_hdmi_in0_frame_cur_word_valid;
assign hdmi2usbsoc_hdmi_in0_frame_frame_valid = hdmi2usbsoc_hdmi_in0_frame_fifo_source_valid;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_source_ready = hdmi2usbsoc_hdmi_in0_frame_frame_ready;
assign hdmi2usbsoc_hdmi_in0_frame_frame_first = hdmi2usbsoc_hdmi_in0_frame_fifo_source_first;
assign hdmi2usbsoc_hdmi_in0_frame_frame_last = hdmi2usbsoc_hdmi_in0_frame_fifo_source_last;
assign hdmi2usbsoc_hdmi_in0_frame_frame_payload_sof = hdmi2usbsoc_hdmi_in0_frame_fifo_source_payload_sof;
assign hdmi2usbsoc_hdmi_in0_frame_frame_payload_pixels = hdmi2usbsoc_hdmi_in0_frame_fifo_source_payload_pixels;
assign hdmi2usbsoc_hdmi_in0_frame_busy = 1'd0;
assign hdmi2usbsoc_hdmi_in0_frame_pix_overflow_reset = hdmi2usbsoc_hdmi_in0_frame_overflow_reset_o;
assign hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_i = hdmi2usbsoc_hdmi_in0_frame_pix_overflow_reset;
assign hdmi2usbsoc_hdmi_in0_frame_overflow_w = (hdmi2usbsoc_hdmi_in0_frame_sys_overflow & (~hdmi2usbsoc_hdmi_in0_frame_overflow_mask));
assign hdmi2usbsoc_hdmi_in0_frame_overflow_reset_i = hdmi2usbsoc_hdmi_in0_frame_overflow_re;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce = (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_ready | (~hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n7));
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_ready = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_valid = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n7;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_busy = ((((((((1'd0 | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n0) | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n1) | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n2) | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n3) | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n4) | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n5) | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n6) | hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n7);
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_first = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n7;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_last = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n7;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_ce = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_r = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_r;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_g = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_g;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_b = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_payload_b;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_y = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_y;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_cb = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cb;
assign hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_payload_cr = hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cr;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce = (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_ready | (~hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n2));
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_ready = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_valid = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n2;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_busy = (((1'd0 | hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n0) | hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n1) | hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n2);
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_first = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n2;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_last = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n2;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_ce = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_y = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_y;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cb = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_cb;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cr = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_payload_cr;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_payload_y = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_y;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_payload_cb_cr = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_cb_cr;
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cb_mean = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cb_sum[8:1];
assign hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cr_mean = hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cr_sum[8:1];
assign hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_din = {hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_last, hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_first, hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_payload_pixels, hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_payload_sof};
assign {hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_last, hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_first, hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_payload_pixels, hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_payload_sof} = hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_dout;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_sink_ready = hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_writable;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_we = hdmi2usbsoc_hdmi_in0_frame_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_first = hdmi2usbsoc_hdmi_in0_frame_fifo_sink_first;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_last = hdmi2usbsoc_hdmi_in0_frame_fifo_sink_last;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_payload_sof = hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_sof;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_in_payload_pixels = hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_pixels;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_source_valid = hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_readable;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_source_first = hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_source_last = hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_source_payload_sof = hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_payload_sof;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_source_payload_pixels = hdmi2usbsoc_hdmi_in0_frame_fifo_fifo_out_payload_pixels;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_re = hdmi2usbsoc_hdmi_in0_frame_fifo_source_ready;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_ce = (hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_writable & hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_we);
assign hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_ce = (hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_readable & hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_re);
assign hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_writable = (((hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q[9] == hdmi2usbsoc_hdmi_in0_frame_fifo_consume_wdomain[9]) | (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q[8] == hdmi2usbsoc_hdmi_in0_frame_fifo_consume_wdomain[8])) | (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q[7:0] != hdmi2usbsoc_hdmi_in0_frame_fifo_consume_wdomain[7:0]));
assign hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_readable = (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q != hdmi2usbsoc_hdmi_in0_frame_fifo_produce_rdomain);
assign hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_adr = hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_binary[8:0];
assign hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_din;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_we = hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_ce;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_rdport_adr = hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary[8:0];
assign hdmi2usbsoc_hdmi_in0_frame_fifo_asyncfifo_dout = hdmi2usbsoc_hdmi_in0_frame_fifo_rdport_dat_r;

// synthesis translate_off
reg dummy_d_87;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next_binary <= 10'd0;
	if (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next_binary <= (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next_binary <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_87 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next = (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next_binary ^ hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_88;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary <= 10'd0;
	if (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary <= (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_88 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next = (hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary ^ hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary[9:1]);
assign hdmi2usbsoc_hdmi_in0_frame_overflow_reset_o = (hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_o ^ hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_o = (hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_o ^ hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_o_r);
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_address_reached = hdmi2usbsoc_hdmi_in0_dma_current_address;
assign hdmi2usbsoc_hdmi_in0_dma_last_word = (hdmi2usbsoc_hdmi_in0_dma_mwords_remaining == 1'd1);
assign hdmi2usbsoc_hdmi_in0_dma_memory_word = {hdmi2usbsoc_hdmi_in0_dma_frame_payload_pixels, hdmi2usbsoc_hdmi_in0_dma_frame_payload_pixels, hdmi2usbsoc_hdmi_in0_dma_frame_payload_pixels, hdmi2usbsoc_hdmi_in0_dma_frame_payload_pixels};
assign hdmi2usbsoc_hdmi_in0_dma_sink_sink_payload_address = hdmi2usbsoc_hdmi_in0_dma_current_address;
assign hdmi2usbsoc_hdmi_in0_dma_sink_sink_payload_data = hdmi2usbsoc_hdmi_in0_dma_memory_word;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_change_slot = ((~hdmi2usbsoc_hdmi_in0_dma_slot_array_address_valid) | hdmi2usbsoc_hdmi_in0_dma_slot_array_address_done);
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_address = comb_rhs_array_muxed36;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_address_valid = comb_rhs_array_muxed37;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_reached = hdmi2usbsoc_hdmi_in0_dma_slot_array_address_reached;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_reached = hdmi2usbsoc_hdmi_in0_dma_slot_array_address_reached;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_done = (hdmi2usbsoc_hdmi_in0_dma_slot_array_address_done & (hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot == 1'd0));
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_done = (hdmi2usbsoc_hdmi_in0_dma_slot_array_address_done & (hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot == 1'd1));

// synthesis translate_off
reg dummy_d_89;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_clear <= 1'd0;
	if ((hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_re & hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_r[0])) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_89 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_90;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_dma_slot_array_status_w <= 2'd0;
	hdmi2usbsoc_hdmi_in0_dma_slot_array_status_w[0] <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status;
	hdmi2usbsoc_hdmi_in0_dma_slot_array_status_w[1] <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status;
// synthesis translate_off
	dummy_d_90 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_91;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_clear <= 1'd0;
	if ((hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_re & hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_r[1])) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_91 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_92;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_w <= 2'd0;
	hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_w[0] <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_pending;
	hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_w[1] <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_pending;
// synthesis translate_off
	dummy_d_92 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_irq = ((hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_w[0] & hdmi2usbsoc_hdmi_in0_dma_slot_array_storage[0]) | (hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_w[1] & hdmi2usbsoc_hdmi_in0_dma_slot_array_storage[1]));
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_trigger;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_pending = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_trigger;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_trigger;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_pending = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_trigger;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_valid = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage[0];
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_dat_w = 2'd2;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_we = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_done;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_dat_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_reached;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_we = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_done;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_trigger = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage[1];
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_valid = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage[0];
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_dat_w = 2'd2;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_we = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_done;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_dat_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_reached;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_we = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_done;
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_trigger = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage[1];
assign hdmi2usbsoc_litedramport0_cmd_payload_we0 = 1'd1;
assign hdmi2usbsoc_litedramport0_cmd_valid0 = (hdmi2usbsoc_hdmi_in0_dma_fifo_sink_ready & hdmi2usbsoc_hdmi_in0_dma_sink_sink_valid);
assign hdmi2usbsoc_litedramport0_cmd_payload_adr0 = hdmi2usbsoc_hdmi_in0_dma_sink_sink_payload_address;
assign hdmi2usbsoc_hdmi_in0_dma_sink_sink_ready = (hdmi2usbsoc_hdmi_in0_dma_fifo_sink_ready & hdmi2usbsoc_litedramport0_cmd_ready0);
assign hdmi2usbsoc_hdmi_in0_dma_fifo_sink_valid = (hdmi2usbsoc_hdmi_in0_dma_sink_sink_valid & hdmi2usbsoc_litedramport0_cmd_ready0);
assign hdmi2usbsoc_hdmi_in0_dma_fifo_sink_payload_data = hdmi2usbsoc_hdmi_in0_dma_sink_sink_payload_data;
assign hdmi2usbsoc_litedramport0_wdata_valid = hdmi2usbsoc_hdmi_in0_dma_fifo_source_valid;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_source_ready = hdmi2usbsoc_litedramport0_wdata_ready;
assign hdmi2usbsoc_litedramport0_wdata_payload_we = 8'd255;
assign hdmi2usbsoc_litedramport0_wdata_payload_data = hdmi2usbsoc_hdmi_in0_dma_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_last, hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_first, hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_last, hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_first, hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_sink_ready = hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_we = hdmi2usbsoc_hdmi_in0_dma_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_first = hdmi2usbsoc_hdmi_in0_dma_fifo_sink_first;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_last = hdmi2usbsoc_hdmi_in0_dma_fifo_sink_last;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_in0_dma_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_source_valid = hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_source_first = hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_source_last = hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_source_payload_data = hdmi2usbsoc_hdmi_in0_dma_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_re = hdmi2usbsoc_hdmi_in0_dma_fifo_source_ready;

// synthesis translate_off
reg dummy_d_93;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_adr <= 4'd0;
	if (hdmi2usbsoc_hdmi_in0_dma_fifo_replace) begin
		hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_in0_dma_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_adr <= hdmi2usbsoc_hdmi_in0_dma_fifo_produce;
	end
// synthesis translate_off
	dummy_d_93 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_we = (hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_in0_dma_fifo_replace));
assign hdmi2usbsoc_hdmi_in0_dma_fifo_do_read = (hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_in0_dma_fifo_rdport_adr = hdmi2usbsoc_hdmi_in0_dma_fifo_consume;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_in0_dma_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_in0_dma_fifo_level != 5'd16);
assign hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_in0_dma_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_94;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in0_dma_reset_words <= 1'd0;
	hdmi2usbsoc_hdmi_in0_dma_count_word <= 1'd0;
	dma0_next_state <= 2'd0;
	hdmi2usbsoc_hdmi_in0_dma_slot_array_address_done <= 1'd0;
	hdmi2usbsoc_hdmi_in0_dma_frame_ready <= 1'd0;
	hdmi2usbsoc_hdmi_in0_dma_sink_sink_valid <= 1'd0;
	dma0_next_state <= dma0_state;
	case (dma0_state)
		1'd1: begin
			hdmi2usbsoc_hdmi_in0_dma_frame_ready <= hdmi2usbsoc_hdmi_in0_dma_sink_sink_ready;
			if (hdmi2usbsoc_hdmi_in0_dma_frame_valid) begin
				hdmi2usbsoc_hdmi_in0_dma_sink_sink_valid <= 1'd1;
				if (hdmi2usbsoc_hdmi_in0_dma_sink_sink_ready) begin
					hdmi2usbsoc_hdmi_in0_dma_count_word <= 1'd1;
					if (hdmi2usbsoc_hdmi_in0_dma_last_word) begin
						dma0_next_state <= 2'd2;
					end
				end
			end
		end
		2'd2: begin
			if ((~hdmi2usbsoc_litedramport0_wdata_valid)) begin
				hdmi2usbsoc_hdmi_in0_dma_slot_array_address_done <= 1'd1;
				dma0_next_state <= 1'd0;
			end
		end
		default: begin
			hdmi2usbsoc_hdmi_in0_dma_reset_words <= 1'd1;
			hdmi2usbsoc_hdmi_in0_dma_frame_ready <= ((~hdmi2usbsoc_hdmi_in0_dma_slot_array_address_valid) | (~hdmi2usbsoc_hdmi_in0_dma_frame_payload_sof));
			if (((hdmi2usbsoc_hdmi_in0_dma_slot_array_address_valid & hdmi2usbsoc_hdmi_in0_dma_frame_payload_sof) & hdmi2usbsoc_hdmi_in0_dma_frame_valid)) begin
				dma0_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_94 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_serdesstrobe = hdmi2usbsoc_hdmi_in1_serdesstrobe;
assign hdmi2usbsoc_hdmi_in1_charsync0_raw_data = hdmi2usbsoc_hdmi_in1_s6datacapture0_d;
assign hdmi2usbsoc_hdmi_in1_wer0_data = hdmi2usbsoc_hdmi_in1_charsync0_data;
assign hdmi2usbsoc_hdmi_in1_decoding0_valid_i = hdmi2usbsoc_hdmi_in1_charsync0_synced;
assign hdmi2usbsoc_hdmi_in1_decoding0_input = hdmi2usbsoc_hdmi_in1_charsync0_data;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_serdesstrobe = hdmi2usbsoc_hdmi_in1_serdesstrobe;
assign hdmi2usbsoc_hdmi_in1_charsync1_raw_data = hdmi2usbsoc_hdmi_in1_s6datacapture1_d;
assign hdmi2usbsoc_hdmi_in1_wer1_data = hdmi2usbsoc_hdmi_in1_charsync1_data;
assign hdmi2usbsoc_hdmi_in1_decoding1_valid_i = hdmi2usbsoc_hdmi_in1_charsync1_synced;
assign hdmi2usbsoc_hdmi_in1_decoding1_input = hdmi2usbsoc_hdmi_in1_charsync1_data;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_serdesstrobe = hdmi2usbsoc_hdmi_in1_serdesstrobe;
assign hdmi2usbsoc_hdmi_in1_charsync2_raw_data = hdmi2usbsoc_hdmi_in1_s6datacapture2_d;
assign hdmi2usbsoc_hdmi_in1_wer2_data = hdmi2usbsoc_hdmi_in1_charsync2_data;
assign hdmi2usbsoc_hdmi_in1_decoding2_valid_i = hdmi2usbsoc_hdmi_in1_charsync2_synced;
assign hdmi2usbsoc_hdmi_in1_decoding2_input = hdmi2usbsoc_hdmi_in1_charsync2_data;
assign hdmi2usbsoc_hdmi_in1_chansync_valid_i = ((hdmi2usbsoc_hdmi_in1_decoding0_valid_o & hdmi2usbsoc_hdmi_in1_decoding1_valid_o) & hdmi2usbsoc_hdmi_in1_decoding2_valid_o);
assign hdmi2usbsoc_hdmi_in1_chansync_data_in0_raw = hdmi2usbsoc_hdmi_in1_decoding0_output_raw;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in0_d = hdmi2usbsoc_hdmi_in1_decoding0_output_d;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in0_c = hdmi2usbsoc_hdmi_in1_decoding0_output_c;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in0_de = hdmi2usbsoc_hdmi_in1_decoding0_output_de;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in1_raw = hdmi2usbsoc_hdmi_in1_decoding1_output_raw;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in1_d = hdmi2usbsoc_hdmi_in1_decoding1_output_d;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in1_c = hdmi2usbsoc_hdmi_in1_decoding1_output_c;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in1_de = hdmi2usbsoc_hdmi_in1_decoding1_output_de;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in2_raw = hdmi2usbsoc_hdmi_in1_decoding2_output_raw;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in2_d = hdmi2usbsoc_hdmi_in1_decoding2_output_d;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in2_c = hdmi2usbsoc_hdmi_in1_decoding2_output_c;
assign hdmi2usbsoc_hdmi_in1_chansync_data_in2_de = hdmi2usbsoc_hdmi_in1_decoding2_output_de;
assign hdmi2usbsoc_hdmi_in1_syncpol_valid_i = hdmi2usbsoc_hdmi_in1_chansync_chan_synced;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in0_raw = hdmi2usbsoc_hdmi_in1_chansync_data_out0_raw;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in0_d = hdmi2usbsoc_hdmi_in1_chansync_data_out0_d;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in0_c = hdmi2usbsoc_hdmi_in1_chansync_data_out0_c;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in0_de = hdmi2usbsoc_hdmi_in1_chansync_data_out0_de;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in1_raw = hdmi2usbsoc_hdmi_in1_chansync_data_out1_raw;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in1_d = hdmi2usbsoc_hdmi_in1_chansync_data_out1_d;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in1_c = hdmi2usbsoc_hdmi_in1_chansync_data_out1_c;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in1_de = hdmi2usbsoc_hdmi_in1_chansync_data_out1_de;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in2_raw = hdmi2usbsoc_hdmi_in1_chansync_data_out2_raw;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in2_d = hdmi2usbsoc_hdmi_in1_chansync_data_out2_d;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in2_c = hdmi2usbsoc_hdmi_in1_chansync_data_out2_c;
assign hdmi2usbsoc_hdmi_in1_syncpol_data_in2_de = hdmi2usbsoc_hdmi_in1_chansync_data_out2_de;
assign hdmi2usbsoc_hdmi_in1_resdetection_valid_i = hdmi2usbsoc_hdmi_in1_syncpol_valid_o;
assign hdmi2usbsoc_hdmi_in1_resdetection_de = hdmi2usbsoc_hdmi_in1_syncpol_de;
assign hdmi2usbsoc_hdmi_in1_resdetection_vsync = hdmi2usbsoc_hdmi_in1_syncpol_vsync;
assign hdmi2usbsoc_hdmi_in1_frame_valid_i = hdmi2usbsoc_hdmi_in1_syncpol_valid_o;
assign hdmi2usbsoc_hdmi_in1_frame_de = hdmi2usbsoc_hdmi_in1_syncpol_de;
assign hdmi2usbsoc_hdmi_in1_frame_vsync = hdmi2usbsoc_hdmi_in1_syncpol_vsync;
assign hdmi2usbsoc_hdmi_in1_frame_r = hdmi2usbsoc_hdmi_in1_syncpol_r;
assign hdmi2usbsoc_hdmi_in1_frame_g = hdmi2usbsoc_hdmi_in1_syncpol_g;
assign hdmi2usbsoc_hdmi_in1_frame_b = hdmi2usbsoc_hdmi_in1_syncpol_b;
assign hdmi2usbsoc_hdmi_in1_dma_frame_valid = hdmi2usbsoc_hdmi_in1_frame_frame_valid;
assign hdmi2usbsoc_hdmi_in1_frame_frame_ready = hdmi2usbsoc_hdmi_in1_dma_frame_ready;
assign hdmi2usbsoc_hdmi_in1_dma_frame_first = hdmi2usbsoc_hdmi_in1_frame_frame_first;
assign hdmi2usbsoc_hdmi_in1_dma_frame_last = hdmi2usbsoc_hdmi_in1_frame_frame_last;
assign hdmi2usbsoc_hdmi_in1_dma_frame_payload_sof = hdmi2usbsoc_hdmi_in1_frame_frame_payload_sof;
assign hdmi2usbsoc_hdmi_in1_dma_frame_payload_pixels = hdmi2usbsoc_hdmi_in1_frame_frame_payload_pixels;
assign hdmi2usbsoc_hdmi_in1_edid_status = 1'd1;
assign hdmi2usbsoc_hdmi_in1_edid_sda_o = (~hdmi2usbsoc_hdmi_in1_edid_sda_drv_reg);
assign hdmi2usbsoc_hdmi_in1_edid_scl_rising = (hdmi2usbsoc_hdmi_in1_edid_scl_i & (~hdmi2usbsoc_hdmi_in1_edid_scl_r));
assign hdmi2usbsoc_hdmi_in1_edid_sda_rising = (hdmi2usbsoc_hdmi_in1_edid_sda_i & (~hdmi2usbsoc_hdmi_in1_edid_sda_r));
assign hdmi2usbsoc_hdmi_in1_edid_sda_falling = ((~hdmi2usbsoc_hdmi_in1_edid_sda_i) & hdmi2usbsoc_hdmi_in1_edid_sda_r);
assign hdmi2usbsoc_hdmi_in1_edid_start = (hdmi2usbsoc_hdmi_in1_edid_scl_i & hdmi2usbsoc_hdmi_in1_edid_sda_falling);
assign hdmi2usbsoc_hdmi_in1_edid_adr = hdmi2usbsoc_hdmi_in1_edid_offset_counter;

// synthesis translate_off
reg dummy_d_95;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_edid_sda_drv <= 1'd0;
	if (hdmi2usbsoc_hdmi_in1_edid_zero_drv) begin
		hdmi2usbsoc_hdmi_in1_edid_sda_drv <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_edid_data_drv) begin
			hdmi2usbsoc_hdmi_in1_edid_sda_drv <= (~hdmi2usbsoc_hdmi_in1_edid_data_bit);
		end
	end
// synthesis translate_off
	dummy_d_95 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_96;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_edid_zero_drv <= 1'd0;
	hdmi2usbsoc_hdmi_in1_edid_data_drv_en <= 1'd0;
	hdmi2usbsoc_hdmi_in1_edid_data_drv_stop <= 1'd0;
	hdmi2usbsoc_hdmi_in1_edid_update_is_read <= 1'd0;
	edid1_next_state <= 4'd0;
	hdmi2usbsoc_hdmi_in1_edid_oc_load <= 1'd0;
	hdmi2usbsoc_hdmi_in1_edid_oc_inc <= 1'd0;
	edid1_next_state <= edid1_state;
	case (edid1_state)
		1'd1: begin
			if ((hdmi2usbsoc_hdmi_in1_edid_counter == 4'd8)) begin
				if ((hdmi2usbsoc_hdmi_in1_edid_din[7:1] == 7'd80)) begin
					hdmi2usbsoc_hdmi_in1_edid_update_is_read <= 1'd1;
					edid1_next_state <= 2'd2;
				end else begin
					edid1_next_state <= 1'd0;
				end
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		2'd2: begin
			if ((~hdmi2usbsoc_hdmi_in1_edid_scl_i)) begin
				edid1_next_state <= 2'd3;
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		2'd3: begin
			hdmi2usbsoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if (hdmi2usbsoc_hdmi_in1_edid_scl_i) begin
				edid1_next_state <= 3'd4;
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		3'd4: begin
			hdmi2usbsoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if ((~hdmi2usbsoc_hdmi_in1_edid_scl_i)) begin
				if (hdmi2usbsoc_hdmi_in1_edid_is_read) begin
					edid1_next_state <= 4'd9;
				end else begin
					edid1_next_state <= 3'd5;
				end
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		3'd5: begin
			if ((hdmi2usbsoc_hdmi_in1_edid_counter == 4'd8)) begin
				hdmi2usbsoc_hdmi_in1_edid_oc_load <= 1'd1;
				edid1_next_state <= 3'd6;
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		3'd6: begin
			if ((~hdmi2usbsoc_hdmi_in1_edid_scl_i)) begin
				edid1_next_state <= 3'd7;
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		3'd7: begin
			hdmi2usbsoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if (hdmi2usbsoc_hdmi_in1_edid_scl_i) begin
				edid1_next_state <= 4'd8;
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		4'd8: begin
			hdmi2usbsoc_hdmi_in1_edid_zero_drv <= 1'd1;
			if ((~hdmi2usbsoc_hdmi_in1_edid_scl_i)) begin
				edid1_next_state <= 1'd1;
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		4'd9: begin
			if ((~hdmi2usbsoc_hdmi_in1_edid_scl_i)) begin
				if ((hdmi2usbsoc_hdmi_in1_edid_counter == 4'd8)) begin
					hdmi2usbsoc_hdmi_in1_edid_data_drv_stop <= 1'd1;
					edid1_next_state <= 4'd10;
				end else begin
					hdmi2usbsoc_hdmi_in1_edid_data_drv_en <= 1'd1;
				end
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		4'd10: begin
			if (hdmi2usbsoc_hdmi_in1_edid_scl_rising) begin
				hdmi2usbsoc_hdmi_in1_edid_oc_inc <= 1'd1;
				if (hdmi2usbsoc_hdmi_in1_edid_sda_i) begin
					edid1_next_state <= 1'd0;
				end else begin
					edid1_next_state <= 4'd9;
				end
			end
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
		default: begin
			if (hdmi2usbsoc_hdmi_in1_edid_start) begin
				edid1_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_96 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_locked_status = hdmi2usbsoc_hdmi_in1_locked;
assign hdmi_in1_pix_o_clk = hdmi_in1_pix_clk;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_too_late = (hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness == 8'd255);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_too_early = (hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness == 1'd0);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_cal = hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_rst = hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_cal = hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_rst = hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_inc = hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_ce = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_o | hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_o);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_i = (hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r[0]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_i = (hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r[1]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_i = (hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r[2]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_i = (hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r[3]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_i = (hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r[4]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_i = (hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r[5]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_busy_status = {hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_slave_pending, hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_master_pending};
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_reset_lateness = hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_i = hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_reset_re;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_o = (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_charsync0_raw = {hdmi2usbsoc_hdmi_in1_charsync0_raw_data, hdmi2usbsoc_hdmi_in1_charsync0_raw_data1};

// synthesis translate_off
reg dummy_d_97;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_wer0_transitions <= 8'd0;
	hdmi2usbsoc_hdmi_in1_wer0_transitions[0] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[0] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[1]);
	hdmi2usbsoc_hdmi_in1_wer0_transitions[1] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[1] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[2]);
	hdmi2usbsoc_hdmi_in1_wer0_transitions[2] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[2] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[3]);
	hdmi2usbsoc_hdmi_in1_wer0_transitions[3] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[3] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[4]);
	hdmi2usbsoc_hdmi_in1_wer0_transitions[4] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[4] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[5]);
	hdmi2usbsoc_hdmi_in1_wer0_transitions[5] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[5] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[6]);
	hdmi2usbsoc_hdmi_in1_wer0_transitions[6] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[6] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[7]);
	hdmi2usbsoc_hdmi_in1_wer0_transitions[7] <= (hdmi2usbsoc_hdmi_in1_wer0_data_r[7] ^ hdmi2usbsoc_hdmi_in1_wer0_data_r[8]);
// synthesis translate_off
	dummy_d_97 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_wer0_i = hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r_updated;
assign hdmi2usbsoc_hdmi_in1_wer0_o = (hdmi2usbsoc_hdmi_in1_wer0_toggle_o ^ hdmi2usbsoc_hdmi_in1_wer0_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_too_late = (hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness == 8'd255);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_too_early = (hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness == 1'd0);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_cal = hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_rst = hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_cal = hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_rst = hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_inc = hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_ce = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_o | hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_o);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_i = (hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r[0]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_i = (hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r[1]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_i = (hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r[2]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_i = (hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r[3]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_i = (hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r[4]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_i = (hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r[5]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_busy_status = {hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_slave_pending, hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_master_pending};
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_reset_lateness = hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_i = hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_reset_re;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_o = (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_charsync1_raw = {hdmi2usbsoc_hdmi_in1_charsync1_raw_data, hdmi2usbsoc_hdmi_in1_charsync1_raw_data1};

// synthesis translate_off
reg dummy_d_98;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_wer1_transitions <= 8'd0;
	hdmi2usbsoc_hdmi_in1_wer1_transitions[0] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[0] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[1]);
	hdmi2usbsoc_hdmi_in1_wer1_transitions[1] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[1] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[2]);
	hdmi2usbsoc_hdmi_in1_wer1_transitions[2] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[2] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[3]);
	hdmi2usbsoc_hdmi_in1_wer1_transitions[3] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[3] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[4]);
	hdmi2usbsoc_hdmi_in1_wer1_transitions[4] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[4] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[5]);
	hdmi2usbsoc_hdmi_in1_wer1_transitions[5] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[5] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[6]);
	hdmi2usbsoc_hdmi_in1_wer1_transitions[6] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[6] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[7]);
	hdmi2usbsoc_hdmi_in1_wer1_transitions[7] <= (hdmi2usbsoc_hdmi_in1_wer1_data_r[7] ^ hdmi2usbsoc_hdmi_in1_wer1_data_r[8]);
// synthesis translate_off
	dummy_d_98 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_wer1_i = hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r_updated;
assign hdmi2usbsoc_hdmi_in1_wer1_o = (hdmi2usbsoc_hdmi_in1_wer1_toggle_o ^ hdmi2usbsoc_hdmi_in1_wer1_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_too_late = (hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness == 8'd255);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_too_early = (hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness == 1'd0);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_cal = hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_rst = hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_cal = hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_rst = hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_inc = hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_ce = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_o | hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_o);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_i = (hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r[0]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_i = (hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r[1]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_i = (hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r[2]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_i = (hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r[3]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_i = (hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r[4]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_i = (hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re & hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r[5]);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_busy_status = {hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_slave_pending, hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_master_pending};
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_reset_lateness = hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_o;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_i = hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_reset_re;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_o = (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_o ^ hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_charsync2_raw = {hdmi2usbsoc_hdmi_in1_charsync2_raw_data, hdmi2usbsoc_hdmi_in1_charsync2_raw_data1};

// synthesis translate_off
reg dummy_d_99;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_wer2_transitions <= 8'd0;
	hdmi2usbsoc_hdmi_in1_wer2_transitions[0] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[0] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[1]);
	hdmi2usbsoc_hdmi_in1_wer2_transitions[1] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[1] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[2]);
	hdmi2usbsoc_hdmi_in1_wer2_transitions[2] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[2] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[3]);
	hdmi2usbsoc_hdmi_in1_wer2_transitions[3] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[3] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[4]);
	hdmi2usbsoc_hdmi_in1_wer2_transitions[4] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[4] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[5]);
	hdmi2usbsoc_hdmi_in1_wer2_transitions[5] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[5] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[6]);
	hdmi2usbsoc_hdmi_in1_wer2_transitions[6] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[6] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[7]);
	hdmi2usbsoc_hdmi_in1_wer2_transitions[7] <= (hdmi2usbsoc_hdmi_in1_wer2_data_r[7] ^ hdmi2usbsoc_hdmi_in1_wer2_data_r[8]);
// synthesis translate_off
	dummy_d_99 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_wer2_i = hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r_updated;
assign hdmi2usbsoc_hdmi_in1_wer2_o = (hdmi2usbsoc_hdmi_in1_wer2_toggle_o ^ hdmi2usbsoc_hdmi_in1_wer2_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_din = {hdmi2usbsoc_hdmi_in1_chansync_data_in0_de, hdmi2usbsoc_hdmi_in1_chansync_data_in0_c, hdmi2usbsoc_hdmi_in1_chansync_data_in0_d, hdmi2usbsoc_hdmi_in1_chansync_data_in0_raw};
assign {hdmi2usbsoc_hdmi_in1_chansync_data_out0_de, hdmi2usbsoc_hdmi_in1_chansync_data_out0_c, hdmi2usbsoc_hdmi_in1_chansync_data_out0_d, hdmi2usbsoc_hdmi_in1_chansync_data_out0_raw} = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_dout;
assign hdmi2usbsoc_hdmi_in1_chansync_is_control0 = (~hdmi2usbsoc_hdmi_in1_chansync_data_out0_de);
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_re = ((~hdmi2usbsoc_hdmi_in1_chansync_is_control0) | hdmi2usbsoc_hdmi_in1_chansync_all_control);
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_din = {hdmi2usbsoc_hdmi_in1_chansync_data_in1_de, hdmi2usbsoc_hdmi_in1_chansync_data_in1_c, hdmi2usbsoc_hdmi_in1_chansync_data_in1_d, hdmi2usbsoc_hdmi_in1_chansync_data_in1_raw};
assign {hdmi2usbsoc_hdmi_in1_chansync_data_out1_de, hdmi2usbsoc_hdmi_in1_chansync_data_out1_c, hdmi2usbsoc_hdmi_in1_chansync_data_out1_d, hdmi2usbsoc_hdmi_in1_chansync_data_out1_raw} = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_dout;
assign hdmi2usbsoc_hdmi_in1_chansync_is_control1 = (~hdmi2usbsoc_hdmi_in1_chansync_data_out1_de);
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_re = ((~hdmi2usbsoc_hdmi_in1_chansync_is_control1) | hdmi2usbsoc_hdmi_in1_chansync_all_control);
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_din = {hdmi2usbsoc_hdmi_in1_chansync_data_in2_de, hdmi2usbsoc_hdmi_in1_chansync_data_in2_c, hdmi2usbsoc_hdmi_in1_chansync_data_in2_d, hdmi2usbsoc_hdmi_in1_chansync_data_in2_raw};
assign {hdmi2usbsoc_hdmi_in1_chansync_data_out2_de, hdmi2usbsoc_hdmi_in1_chansync_data_out2_c, hdmi2usbsoc_hdmi_in1_chansync_data_out2_d, hdmi2usbsoc_hdmi_in1_chansync_data_out2_raw} = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_dout;
assign hdmi2usbsoc_hdmi_in1_chansync_is_control2 = (~hdmi2usbsoc_hdmi_in1_chansync_data_out2_de);
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_re = ((~hdmi2usbsoc_hdmi_in1_chansync_is_control2) | hdmi2usbsoc_hdmi_in1_chansync_all_control);
assign hdmi2usbsoc_hdmi_in1_chansync_all_control = ((hdmi2usbsoc_hdmi_in1_chansync_is_control0 & hdmi2usbsoc_hdmi_in1_chansync_is_control1) & hdmi2usbsoc_hdmi_in1_chansync_is_control2);
assign hdmi2usbsoc_hdmi_in1_chansync_some_control = ((hdmi2usbsoc_hdmi_in1_chansync_is_control0 | hdmi2usbsoc_hdmi_in1_chansync_is_control1) | hdmi2usbsoc_hdmi_in1_chansync_is_control2);
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_adr = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_produce;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_w = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_din;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_we = 1'd1;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_rdport_adr = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_consume;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_dout = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_adr = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_produce;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_w = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_din;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_we = 1'd1;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_rdport_adr = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_consume;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_dout = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_adr = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_produce;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_w = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_din;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_we = 1'd1;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_rdport_adr = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_consume;
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_dout = hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in1_syncpol_de = hdmi2usbsoc_hdmi_in1_syncpol_de_r;
assign hdmi2usbsoc_hdmi_in1_syncpol_hsync = hdmi2usbsoc_hdmi_in1_syncpol_c_out[0];
assign hdmi2usbsoc_hdmi_in1_syncpol_vsync = hdmi2usbsoc_hdmi_in1_syncpol_c_out[1];
assign hdmi2usbsoc_hdmi_in1_resdetection_pn_de = ((~hdmi2usbsoc_hdmi_in1_resdetection_de) & hdmi2usbsoc_hdmi_in1_resdetection_de_r);
assign hdmi2usbsoc_hdmi_in1_resdetection_p_vsync = (hdmi2usbsoc_hdmi_in1_resdetection_vsync & (~hdmi2usbsoc_hdmi_in1_resdetection_vsync_r));
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_valid = hdmi2usbsoc_hdmi_in1_frame_valid_i;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_r = hdmi2usbsoc_hdmi_in1_frame_r;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_g = hdmi2usbsoc_hdmi_in1_frame_g;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_b = hdmi2usbsoc_hdmi_in1_frame_b;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_valid = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_valid;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_ready = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_ready;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_first = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_first;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_last = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_last;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_y = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_y;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_cb = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_cb;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_cr = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_cr;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_ready = 1'd1;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first = (hdmi2usbsoc_hdmi_in1_frame_de & (~hdmi2usbsoc_hdmi_in1_frame_de_r));
assign hdmi2usbsoc_hdmi_in1_frame_new_frame = (hdmi2usbsoc_hdmi_in1_frame_next_vsync10 & (~hdmi2usbsoc_hdmi_in1_frame_vsync_r));
assign hdmi2usbsoc_hdmi_in1_frame_encoded_pixel = {hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_payload_cb_cr, hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_payload_y};
assign hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_pixels = hdmi2usbsoc_hdmi_in1_frame_cur_word;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_sink_valid = hdmi2usbsoc_hdmi_in1_frame_cur_word_valid;
assign hdmi2usbsoc_hdmi_in1_frame_frame_valid = hdmi2usbsoc_hdmi_in1_frame_fifo_source_valid;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_source_ready = hdmi2usbsoc_hdmi_in1_frame_frame_ready;
assign hdmi2usbsoc_hdmi_in1_frame_frame_first = hdmi2usbsoc_hdmi_in1_frame_fifo_source_first;
assign hdmi2usbsoc_hdmi_in1_frame_frame_last = hdmi2usbsoc_hdmi_in1_frame_fifo_source_last;
assign hdmi2usbsoc_hdmi_in1_frame_frame_payload_sof = hdmi2usbsoc_hdmi_in1_frame_fifo_source_payload_sof;
assign hdmi2usbsoc_hdmi_in1_frame_frame_payload_pixels = hdmi2usbsoc_hdmi_in1_frame_fifo_source_payload_pixels;
assign hdmi2usbsoc_hdmi_in1_frame_busy = 1'd0;
assign hdmi2usbsoc_hdmi_in1_frame_pix_overflow_reset = hdmi2usbsoc_hdmi_in1_frame_overflow_reset_o;
assign hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_i = hdmi2usbsoc_hdmi_in1_frame_pix_overflow_reset;
assign hdmi2usbsoc_hdmi_in1_frame_overflow_w = (hdmi2usbsoc_hdmi_in1_frame_sys_overflow & (~hdmi2usbsoc_hdmi_in1_frame_overflow_mask));
assign hdmi2usbsoc_hdmi_in1_frame_overflow_reset_i = hdmi2usbsoc_hdmi_in1_frame_overflow_re;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce = (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_ready | (~hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n7));
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_ready = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_valid = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n7;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_busy = ((((((((1'd0 | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n0) | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n1) | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n2) | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n3) | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n4) | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n5) | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n6) | hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n7);
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_first = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n7;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_last = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n7;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_ce = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_r = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_r;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_g = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_g;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_b = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_payload_b;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_y = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_y;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_cb = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cb;
assign hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_payload_cr = hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cr;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce = (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_ready | (~hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n2));
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_ready = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_valid = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n2;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_busy = (((1'd0 | hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n0) | hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n1) | hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n2);
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_first = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n2;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_last = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n2;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_ce = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_y = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_y;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cb = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_cb;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cr = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_payload_cr;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_payload_y = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_y;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_payload_cb_cr = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_cb_cr;
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cb_mean = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cb_sum[8:1];
assign hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cr_mean = hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cr_sum[8:1];
assign hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_din = {hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_last, hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_first, hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_payload_pixels, hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_payload_sof};
assign {hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_last, hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_first, hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_payload_pixels, hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_payload_sof} = hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_dout;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_sink_ready = hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_writable;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_we = hdmi2usbsoc_hdmi_in1_frame_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_first = hdmi2usbsoc_hdmi_in1_frame_fifo_sink_first;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_last = hdmi2usbsoc_hdmi_in1_frame_fifo_sink_last;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_payload_sof = hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_sof;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_in_payload_pixels = hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_pixels;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_source_valid = hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_readable;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_source_first = hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_source_last = hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_source_payload_sof = hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_payload_sof;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_source_payload_pixels = hdmi2usbsoc_hdmi_in1_frame_fifo_fifo_out_payload_pixels;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_re = hdmi2usbsoc_hdmi_in1_frame_fifo_source_ready;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_ce = (hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_writable & hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_we);
assign hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_ce = (hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_readable & hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_re);
assign hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_writable = (((hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q[9] == hdmi2usbsoc_hdmi_in1_frame_fifo_consume_wdomain[9]) | (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q[8] == hdmi2usbsoc_hdmi_in1_frame_fifo_consume_wdomain[8])) | (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q[7:0] != hdmi2usbsoc_hdmi_in1_frame_fifo_consume_wdomain[7:0]));
assign hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_readable = (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q != hdmi2usbsoc_hdmi_in1_frame_fifo_produce_rdomain);
assign hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_adr = hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_binary[8:0];
assign hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_din;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_we = hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_ce;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_rdport_adr = hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary[8:0];
assign hdmi2usbsoc_hdmi_in1_frame_fifo_asyncfifo_dout = hdmi2usbsoc_hdmi_in1_frame_fifo_rdport_dat_r;

// synthesis translate_off
reg dummy_d_100;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next_binary <= 10'd0;
	if (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next_binary <= (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next_binary <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_100 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next = (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next_binary ^ hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_101;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary <= 10'd0;
	if (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary <= (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_101 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next = (hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary ^ hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary[9:1]);
assign hdmi2usbsoc_hdmi_in1_frame_overflow_reset_o = (hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_o ^ hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_o = (hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_o ^ hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_o_r);
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_address_reached = hdmi2usbsoc_hdmi_in1_dma_current_address;
assign hdmi2usbsoc_hdmi_in1_dma_last_word = (hdmi2usbsoc_hdmi_in1_dma_mwords_remaining == 1'd1);
assign hdmi2usbsoc_hdmi_in1_dma_memory_word = {hdmi2usbsoc_hdmi_in1_dma_frame_payload_pixels, hdmi2usbsoc_hdmi_in1_dma_frame_payload_pixels, hdmi2usbsoc_hdmi_in1_dma_frame_payload_pixels, hdmi2usbsoc_hdmi_in1_dma_frame_payload_pixels};
assign hdmi2usbsoc_hdmi_in1_dma_sink_sink_payload_address = hdmi2usbsoc_hdmi_in1_dma_current_address;
assign hdmi2usbsoc_hdmi_in1_dma_sink_sink_payload_data = hdmi2usbsoc_hdmi_in1_dma_memory_word;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_change_slot = ((~hdmi2usbsoc_hdmi_in1_dma_slot_array_address_valid) | hdmi2usbsoc_hdmi_in1_dma_slot_array_address_done);
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_address = comb_rhs_array_muxed38;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_address_valid = comb_rhs_array_muxed39;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_reached = hdmi2usbsoc_hdmi_in1_dma_slot_array_address_reached;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_reached = hdmi2usbsoc_hdmi_in1_dma_slot_array_address_reached;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_done = (hdmi2usbsoc_hdmi_in1_dma_slot_array_address_done & (hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot == 1'd0));
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_done = (hdmi2usbsoc_hdmi_in1_dma_slot_array_address_done & (hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot == 1'd1));

// synthesis translate_off
reg dummy_d_102;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_clear <= 1'd0;
	if ((hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_re & hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_r[0])) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_102 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_103;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_dma_slot_array_status_w <= 2'd0;
	hdmi2usbsoc_hdmi_in1_dma_slot_array_status_w[0] <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status;
	hdmi2usbsoc_hdmi_in1_dma_slot_array_status_w[1] <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status;
// synthesis translate_off
	dummy_d_103 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_104;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_clear <= 1'd0;
	if ((hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_re & hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_r[1])) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_104 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_105;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_w <= 2'd0;
	hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_w[0] <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_pending;
	hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_w[1] <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_pending;
// synthesis translate_off
	dummy_d_105 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_irq = ((hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_w[0] & hdmi2usbsoc_hdmi_in1_dma_slot_array_storage[0]) | (hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_w[1] & hdmi2usbsoc_hdmi_in1_dma_slot_array_storage[1]));
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_trigger;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_pending = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_trigger;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_trigger;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_pending = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_trigger;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_valid = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage[0];
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_dat_w = 2'd2;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_we = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_done;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_dat_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_reached;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_we = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_done;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_trigger = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage[1];
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_valid = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage[0];
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_dat_w = 2'd2;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_we = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_done;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_dat_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_reached;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_we = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_done;
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_trigger = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage[1];
assign hdmi2usbsoc_litedramport1_cmd_payload_we0 = 1'd1;
assign hdmi2usbsoc_litedramport1_cmd_valid0 = (hdmi2usbsoc_hdmi_in1_dma_fifo_sink_ready & hdmi2usbsoc_hdmi_in1_dma_sink_sink_valid);
assign hdmi2usbsoc_litedramport1_cmd_payload_adr0 = hdmi2usbsoc_hdmi_in1_dma_sink_sink_payload_address;
assign hdmi2usbsoc_hdmi_in1_dma_sink_sink_ready = (hdmi2usbsoc_hdmi_in1_dma_fifo_sink_ready & hdmi2usbsoc_litedramport1_cmd_ready0);
assign hdmi2usbsoc_hdmi_in1_dma_fifo_sink_valid = (hdmi2usbsoc_hdmi_in1_dma_sink_sink_valid & hdmi2usbsoc_litedramport1_cmd_ready0);
assign hdmi2usbsoc_hdmi_in1_dma_fifo_sink_payload_data = hdmi2usbsoc_hdmi_in1_dma_sink_sink_payload_data;
assign hdmi2usbsoc_litedramport1_wdata_valid = hdmi2usbsoc_hdmi_in1_dma_fifo_source_valid;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_source_ready = hdmi2usbsoc_litedramport1_wdata_ready;
assign hdmi2usbsoc_litedramport1_wdata_payload_we = 8'd255;
assign hdmi2usbsoc_litedramport1_wdata_payload_data = hdmi2usbsoc_hdmi_in1_dma_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_last, hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_first, hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_last, hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_first, hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_sink_ready = hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_we = hdmi2usbsoc_hdmi_in1_dma_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_first = hdmi2usbsoc_hdmi_in1_dma_fifo_sink_first;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_last = hdmi2usbsoc_hdmi_in1_dma_fifo_sink_last;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_in1_dma_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_source_valid = hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_source_first = hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_source_last = hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_source_payload_data = hdmi2usbsoc_hdmi_in1_dma_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_re = hdmi2usbsoc_hdmi_in1_dma_fifo_source_ready;

// synthesis translate_off
reg dummy_d_106;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_adr <= 4'd0;
	if (hdmi2usbsoc_hdmi_in1_dma_fifo_replace) begin
		hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_in1_dma_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_adr <= hdmi2usbsoc_hdmi_in1_dma_fifo_produce;
	end
// synthesis translate_off
	dummy_d_106 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_we = (hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_in1_dma_fifo_replace));
assign hdmi2usbsoc_hdmi_in1_dma_fifo_do_read = (hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_in1_dma_fifo_rdport_adr = hdmi2usbsoc_hdmi_in1_dma_fifo_consume;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_in1_dma_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_in1_dma_fifo_level != 5'd16);
assign hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_in1_dma_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_107;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_in1_dma_sink_sink_valid <= 1'd0;
	dma1_next_state <= 2'd0;
	hdmi2usbsoc_hdmi_in1_dma_reset_words <= 1'd0;
	hdmi2usbsoc_hdmi_in1_dma_count_word <= 1'd0;
	hdmi2usbsoc_hdmi_in1_dma_slot_array_address_done <= 1'd0;
	hdmi2usbsoc_hdmi_in1_dma_frame_ready <= 1'd0;
	dma1_next_state <= dma1_state;
	case (dma1_state)
		1'd1: begin
			hdmi2usbsoc_hdmi_in1_dma_frame_ready <= hdmi2usbsoc_hdmi_in1_dma_sink_sink_ready;
			if (hdmi2usbsoc_hdmi_in1_dma_frame_valid) begin
				hdmi2usbsoc_hdmi_in1_dma_sink_sink_valid <= 1'd1;
				if (hdmi2usbsoc_hdmi_in1_dma_sink_sink_ready) begin
					hdmi2usbsoc_hdmi_in1_dma_count_word <= 1'd1;
					if (hdmi2usbsoc_hdmi_in1_dma_last_word) begin
						dma1_next_state <= 2'd2;
					end
				end
			end
		end
		2'd2: begin
			if ((~hdmi2usbsoc_litedramport1_wdata_valid)) begin
				hdmi2usbsoc_hdmi_in1_dma_slot_array_address_done <= 1'd1;
				dma1_next_state <= 1'd0;
			end
		end
		default: begin
			hdmi2usbsoc_hdmi_in1_dma_reset_words <= 1'd1;
			hdmi2usbsoc_hdmi_in1_dma_frame_ready <= ((~hdmi2usbsoc_hdmi_in1_dma_slot_array_address_valid) | (~hdmi2usbsoc_hdmi_in1_dma_frame_payload_sof));
			if (((hdmi2usbsoc_hdmi_in1_dma_slot_array_address_valid & hdmi2usbsoc_hdmi_in1_dma_frame_payload_sof) & hdmi2usbsoc_hdmi_in1_dma_frame_valid)) begin
				dma1_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_107 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_core_source_source_ready = 1'd1;
assign hdmi2usbsoc_hdmi_out0_resetinserter_reset = (hdmi2usbsoc_hdmi_out0_core_source_source_param_de & (~hdmi2usbsoc_hdmi_out0_de_r));
assign hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_valid = hdmi2usbsoc_hdmi_out0_core_source_valid_d;
assign hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_y = hdmi2usbsoc_hdmi_out0_core_source_data_d[7:0];
assign hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr = hdmi2usbsoc_hdmi_out0_core_source_data_d[15:8];
assign hdmi2usbsoc_hdmi_out0_sink_valid = hdmi2usbsoc_hdmi_out0_resetinserter_source_source_valid;
assign hdmi2usbsoc_hdmi_out0_resetinserter_source_source_ready = hdmi2usbsoc_hdmi_out0_sink_ready;
assign hdmi2usbsoc_hdmi_out0_sink_first = hdmi2usbsoc_hdmi_out0_resetinserter_source_source_first;
assign hdmi2usbsoc_hdmi_out0_sink_last = hdmi2usbsoc_hdmi_out0_resetinserter_source_source_last;
assign hdmi2usbsoc_hdmi_out0_sink_payload_y = hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_y;
assign hdmi2usbsoc_hdmi_out0_sink_payload_cb = hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_cb;
assign hdmi2usbsoc_hdmi_out0_sink_payload_cr = hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_cr;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_valid = hdmi2usbsoc_hdmi_out0_source_valid;
assign hdmi2usbsoc_hdmi_out0_source_ready = hdmi2usbsoc_hdmi_out0_driver_sink_sink_ready;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_first = hdmi2usbsoc_hdmi_out0_source_first;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_last = hdmi2usbsoc_hdmi_out0_source_last;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_r = hdmi2usbsoc_hdmi_out0_source_payload_r;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_g = hdmi2usbsoc_hdmi_out0_source_payload_g;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_b = hdmi2usbsoc_hdmi_out0_source_payload_b;
assign hdmi2usbsoc_hdmi_out0_sink_payload_de = hdmi2usbsoc_hdmi_out0_core_source_source_param_de;
assign hdmi2usbsoc_hdmi_out0_sink_payload_vsync = hdmi2usbsoc_hdmi_out0_core_source_source_param_vsync;
assign hdmi2usbsoc_hdmi_out0_sink_payload_hsync = hdmi2usbsoc_hdmi_out0_core_source_source_param_hsync;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_de = hdmi2usbsoc_hdmi_out0_source_payload_de;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_vsync = hdmi2usbsoc_hdmi_out0_source_payload_vsync;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_hsync = hdmi2usbsoc_hdmi_out0_source_payload_hsync;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_valid = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_valid;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_sink_valid = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_valid;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_ready = hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_ready;
assign hdmi2usbsoc_hdmi_out0_core_source_source_valid = (hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_valid & ((~hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_de) | hdmi2usbsoc_hdmi_out0_core_dmareader_source_valid));

// synthesis translate_off
reg dummy_d_108;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_ready <= 1'd0;
	hdmi2usbsoc_hdmi_out0_core_dmareader_source_ready <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_out0_core_initiator_source_source_valid)) begin
		hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_ready <= 1'd1;
		hdmi2usbsoc_hdmi_out0_core_dmareader_source_ready <= 1'd1;
	end else begin
		if ((hdmi2usbsoc_hdmi_out0_core_source_source_valid & hdmi2usbsoc_hdmi_out0_core_source_source_ready)) begin
			hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_ready <= 1'd1;
			hdmi2usbsoc_hdmi_out0_core_dmareader_source_ready <= (hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_de | 1'd0);
		end
	end
// synthesis translate_off
	dummy_d_108 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hres = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hres;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hscan = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hscan;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vres = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vres;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vscan = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vscan;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_sink_payload_base = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_base;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_sink_payload_length = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_length;
assign hdmi2usbsoc_hdmi_out0_core_source_source_param_de = hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_de;
assign hdmi2usbsoc_hdmi_out0_core_source_source_param_hsync = hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_hsync;
assign hdmi2usbsoc_hdmi_out0_core_source_source_param_vsync = hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_vsync;
assign hdmi2usbsoc_hdmi_out0_core_source_source_payload_data = hdmi2usbsoc_hdmi_out0_core_dmareader_source_payload_data;
assign hdmi2usbsoc_hdmi_out0_core_i = hdmi2usbsoc_hdmi_out0_core_underflow_update_underflow_update_re;
assign hdmi2usbsoc_hdmi_out0_core_underflow_update = hdmi2usbsoc_hdmi_out0_core_o;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hres = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hscan = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vres = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vscan = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_base = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_length = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_valid = hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_valid = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_valid;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_ready = hdmi2usbsoc_hdmi_out0_core_initiator_source_source_ready;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_first = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_first;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_last = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_last;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hres = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hres;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_hscan = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hscan;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vres = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vres;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_vscan = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vscan;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_base = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_base;
assign hdmi2usbsoc_hdmi_out0_core_initiator_source_source_payload_length = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_length;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_din = {hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_last, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_first, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_length, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_base, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vres, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hres};
assign {hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_last, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_first, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_length, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_base, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vres, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start, hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hres} = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_dout;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_ready = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_writable;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_we = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_valid;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_first = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_first;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_last = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_last;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hres = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hres;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_hscan;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vres = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vres;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_vscan;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_base = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_base;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_in_payload_length = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_sink_payload_length;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_valid = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_readable;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_first = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_first;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_last = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_last;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hres = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hres;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_hscan = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vres = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vres;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vsync_start = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vsync_end = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_vscan = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_base = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_base;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_payload_length = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_fifo_out_payload_length;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_re = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_source_ready;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_ce = (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_writable & hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_we);
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_ce = (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_readable & hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_re);
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_writable = ((hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q[1] == hdmi2usbsoc_hdmi_out0_core_initiator_cdc_consume_wdomain[1]) | (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q[0] == hdmi2usbsoc_hdmi_out0_core_initiator_cdc_consume_wdomain[0]));
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_readable = (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q != hdmi2usbsoc_hdmi_out0_core_initiator_cdc_produce_rdomain);
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_adr = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary[0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_dat_w = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_din;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_we = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_ce;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_rdport_adr = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary[0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_asyncfifo_dout = hdmi2usbsoc_hdmi_out0_core_initiator_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_109;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= 2'd0;
	if (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_ce) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_109 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next = (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary ^ hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary[1]);

// synthesis translate_off
reg dummy_d_110;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= 2'd0;
	if (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_ce) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_110 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next = (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary ^ hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary[1]);

// synthesis translate_off
reg dummy_d_111;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_de <= 1'd0;
	hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_valid <= 1'd0;
	hdmi2usbsoc_hdmi_out0_core_timinggenerator_active <= 1'd0;
	if (hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_valid) begin
		hdmi2usbsoc_hdmi_out0_core_timinggenerator_active <= (hdmi2usbsoc_hdmi_out0_core_timinggenerator_hactive & hdmi2usbsoc_hdmi_out0_core_timinggenerator_vactive);
		hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_valid <= 1'd1;
		if (hdmi2usbsoc_hdmi_out0_core_timinggenerator_active) begin
			hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_de <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_111 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_ready = (hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_ready & hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_last);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_base = hdmi2usbsoc_hdmi_out0_core_dmareader_sink_payload_base[31:1];
assign hdmi2usbsoc_hdmi_out0_core_dmareader_length = hdmi2usbsoc_hdmi_out0_core_dmareader_sink_payload_length[31:1];
assign hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_payload_address = (hdmi2usbsoc_hdmi_out0_core_dmareader_base + hdmi2usbsoc_hdmi_out0_core_dmareader_offset);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_valid = hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_valid;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_ready = hdmi2usbsoc_hdmi_out0_core_dmareader_source_ready;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_first = hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_first;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_last = hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_last;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_payload_data = hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_payload_data;
assign hdmi2usbsoc_litedramport1_cmd_payload_we1 = 1'd0;
assign hdmi2usbsoc_litedramport1_cmd_valid1 = (hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_valid & hdmi2usbsoc_hdmi_out0_core_dmareader_request_enable);
assign hdmi2usbsoc_litedramport1_cmd_payload_adr1 = hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_payload_address;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_ready = (hdmi2usbsoc_litedramport1_cmd_ready1 & hdmi2usbsoc_hdmi_out0_core_dmareader_request_enable);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_request_issued = (hdmi2usbsoc_litedramport1_cmd_valid1 & hdmi2usbsoc_litedramport1_cmd_ready1);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_request_enable = (hdmi2usbsoc_hdmi_out0_core_dmareader_rsv_level != 13'd4096);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_valid = hdmi2usbsoc_litedramport1_rdata_valid1;
assign hdmi2usbsoc_litedramport1_rdata_ready = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_ready;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_first = hdmi2usbsoc_litedramport1_rdata_first;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_last = hdmi2usbsoc_litedramport1_rdata_last;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_payload_data = hdmi2usbsoc_litedramport1_rdata_payload_data1;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_valid = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_valid;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_ready = hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_ready;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_first = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_first;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_last = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_last;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_payload_data = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_data_dequeued = (hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_valid & hdmi2usbsoc_hdmi_out0_core_dmareader_source_source_ready);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_ready = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_valid = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_readable;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_first = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_last = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_payload_data = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_re = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_source_ready;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_re = (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_readable & ((~hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_readable) | hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_re));
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level1 = (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 + hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_readable);

// synthesis translate_off
reg dummy_d_112;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_adr <= 12'd0;
	if (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_replace) begin
		hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_produce;
	end
// synthesis translate_off
	dummy_d_112 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_we = (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_replace));
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_do_read = (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_adr = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_consume;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_re = hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_do_read;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 != 13'd4096);
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 != 1'd0);

// synthesis translate_off
reg dummy_d_113;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value_ce <= 1'd0;
	hdmi2usbsoc_hdmi_out0_core_dmareader_sink_ready <= 1'd0;
	hdmi2usbsoc_litedramport1_flush <= 1'd0;
	hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_valid <= 1'd0;
	videoout0_next_state <= 1'd0;
	hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value <= 26'd0;
	videoout0_next_state <= videoout0_state;
	case (videoout0_state)
		1'd1: begin
			hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_valid <= 1'd1;
			if (hdmi2usbsoc_hdmi_out0_core_dmareader_sink_sink_ready) begin
				hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value <= (hdmi2usbsoc_hdmi_out0_core_dmareader_offset + 1'd1);
				hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value_ce <= 1'd1;
				if ((hdmi2usbsoc_hdmi_out0_core_dmareader_offset == (hdmi2usbsoc_hdmi_out0_core_dmareader_length - 1'd1))) begin
					hdmi2usbsoc_hdmi_out0_core_dmareader_sink_ready <= 1'd1;
					videoout0_next_state <= 1'd0;
				end
			end
		end
		default: begin
			hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value <= 1'd0;
			hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value_ce <= 1'd1;
			if (hdmi2usbsoc_hdmi_out0_core_dmareader_sink_valid) begin
				videoout0_next_state <= 1'd1;
			end else begin
				hdmi2usbsoc_litedramport1_flush <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_113 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_core_o = (hdmi2usbsoc_hdmi_out0_core_toggle_o ^ hdmi2usbsoc_hdmi_out0_core_toggle_o_r);
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe = hdmi2usbsoc_hdmi_out0_driver_clocking_serdesstrobe;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_valid = hdmi2usbsoc_hdmi_out0_driver_sink_sink_valid;
assign hdmi2usbsoc_hdmi_out0_driver_sink_sink_ready = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_ready;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_first = hdmi2usbsoc_hdmi_out0_driver_sink_sink_first;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_last = hdmi2usbsoc_hdmi_out0_driver_sink_sink_last;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_r = hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_r;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_g = hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_g;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_b = hdmi2usbsoc_hdmi_out0_driver_sink_sink_payload_b;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_hsync = hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_hsync;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_vsync = hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_vsync;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_de = hdmi2usbsoc_hdmi_out0_driver_sink_sink_param_de;
assign hdmi2usbsoc_hdmi_out0_driver_clocking_transmitting = (hdmi2usbsoc_hdmi_out0_driver_clocking_remaining_bits != 1'd0);
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progdata = (hdmi2usbsoc_hdmi_out0_driver_clocking_transmitting & hdmi2usbsoc_hdmi_out0_driver_clocking_sr[0]);
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progen = (hdmi2usbsoc_hdmi_out0_driver_clocking_transmitting | hdmi2usbsoc_hdmi_out0_driver_clocking_send_go_re);
assign hdmi2usbsoc_hdmi_out0_driver_clocking_busy = (hdmi2usbsoc_hdmi_out0_driver_clocking_busy_counter != 1'd0);
assign hdmi2usbsoc_hdmi_out0_driver_clocking_status_status = {hdmi2usbsoc_hdmi_out0_driver_clocking_mult_locked, hdmi2usbsoc_hdmi_out0_driver_clocking_pix_locked, hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progdone, hdmi2usbsoc_hdmi_out0_driver_clocking_busy};
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_ready = 1'd1;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0 = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_b;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0 = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_g;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0 = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_payload_r;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_c = {hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_vsync, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_hsync};
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_c = 1'd0;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_c = 1'd0;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_de = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_de;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_de = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_de;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_de = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_sink_param_de;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x_pol;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n = ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1d > 3'd4) | ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1d == 3'd4) & (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0])));
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x_pol;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n = ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1d > 3'd4) | ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1d == 3'd4) & (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0])));
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x = hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x_pol;
assign hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n = ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1d > 3'd4) | ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1d == 3'd4) & (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0])));

// synthesis translate_off
reg dummy_d_114;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_valid <= 1'd0;
	hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_valid <= 1'd0;
	hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_valid <= 1'd0;
	hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_payload_data <= 8'd0;
	hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready <= 1'd0;
	hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data <= 8'd0;
	hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data <= 8'd0;
	if ((~hdmi2usbsoc_hdmi_out0_resetinserter_parity_in)) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_y;
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
		hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready <= (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_ready & hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_ready);
	end else begin
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_y;
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
		hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready <= (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_ready & hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_ready);
	end
// synthesis translate_off
	dummy_d_114 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_resetinserter_source_source_valid = ((hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_valid & hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_valid) & hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_valid);
assign hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_y = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_cb = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_source_source_payload_cr = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_ready = (hdmi2usbsoc_hdmi_out0_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out0_resetinserter_source_source_ready);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_ready = ((hdmi2usbsoc_hdmi_out0_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out0_resetinserter_source_source_ready) & hdmi2usbsoc_hdmi_out0_resetinserter_parity_out);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_ready = ((hdmi2usbsoc_hdmi_out0_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out0_resetinserter_source_source_ready) & hdmi2usbsoc_hdmi_out0_resetinserter_parity_out);
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_ready = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_valid = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_first = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_last = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_payload_data = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_re = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_source_ready;

// synthesis translate_off
reg dummy_d_115;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_replace) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_produce;
	end
// synthesis translate_off
	dummy_d_115 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_we = (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_replace));
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_do_read = (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_rdport_adr = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_consume;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level != 3'd4);
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_ready = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_valid = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_first = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_last = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_payload_data = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_re = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_source_ready;

// synthesis translate_off
reg dummy_d_116;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_replace) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_produce;
	end
// synthesis translate_off
	dummy_d_116 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_we = (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_replace));
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_do_read = (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_rdport_adr = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_consume;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level != 3'd4);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_ready = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_valid = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_first = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_last = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_payload_data = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_re = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_source_ready;

// synthesis translate_off
reg dummy_d_117;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_replace) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_produce;
	end
// synthesis translate_off
	dummy_d_117 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_we = (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_replace));
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_do_read = (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_rdport_adr = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_consume;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level != 3'd4);
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi_out0_pipe_ce = (hdmi2usbsoc_hdmi_out0_source_ready | (~hdmi2usbsoc_hdmi_out0_valid_n3));
assign hdmi2usbsoc_hdmi_out0_sink_ready = hdmi2usbsoc_hdmi_out0_pipe_ce;
assign hdmi2usbsoc_hdmi_out0_source_valid = hdmi2usbsoc_hdmi_out0_valid_n3;
assign hdmi2usbsoc_hdmi_out0_busy = ((((1'd0 | hdmi2usbsoc_hdmi_out0_valid_n0) | hdmi2usbsoc_hdmi_out0_valid_n1) | hdmi2usbsoc_hdmi_out0_valid_n2) | hdmi2usbsoc_hdmi_out0_valid_n3);
assign hdmi2usbsoc_hdmi_out0_source_first = hdmi2usbsoc_hdmi_out0_first_n3;
assign hdmi2usbsoc_hdmi_out0_source_last = hdmi2usbsoc_hdmi_out0_last_n3;
assign hdmi2usbsoc_hdmi_out0_ce = hdmi2usbsoc_hdmi_out0_pipe_ce;
assign hdmi2usbsoc_hdmi_out0_sink_y = hdmi2usbsoc_hdmi_out0_sink_payload_y;
assign hdmi2usbsoc_hdmi_out0_sink_cb = hdmi2usbsoc_hdmi_out0_sink_payload_cb;
assign hdmi2usbsoc_hdmi_out0_sink_cr = hdmi2usbsoc_hdmi_out0_sink_payload_cr;
assign hdmi2usbsoc_hdmi_out0_source_payload_r = hdmi2usbsoc_hdmi_out0_source_r;
assign hdmi2usbsoc_hdmi_out0_source_payload_g = hdmi2usbsoc_hdmi_out0_source_g;
assign hdmi2usbsoc_hdmi_out0_source_payload_b = hdmi2usbsoc_hdmi_out0_source_b;
assign hdmi2usbsoc_hdmi_out0_source_payload_hsync = hdmi2usbsoc_hdmi_out0_next_s5;
assign hdmi2usbsoc_hdmi_out0_source_payload_vsync = hdmi2usbsoc_hdmi_out0_next_s11;
assign hdmi2usbsoc_hdmi_out0_source_payload_de = hdmi2usbsoc_hdmi_out0_next_s17;
assign hdmi2usbsoc_hdmi_out1_core_source_source_ready = 1'd1;
assign hdmi2usbsoc_hdmi_out1_resetinserter_reset = (hdmi2usbsoc_hdmi_out1_core_source_source_param_de & (~hdmi2usbsoc_hdmi_out1_de_r));
assign hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_valid = hdmi2usbsoc_hdmi_out1_core_source_valid_d;
assign hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_y = hdmi2usbsoc_hdmi_out1_core_source_data_d[7:0];
assign hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_cb_cr = hdmi2usbsoc_hdmi_out1_core_source_data_d[15:8];
assign hdmi2usbsoc_hdmi_out1_sink_valid = hdmi2usbsoc_hdmi_out1_resetinserter_source_source_valid;
assign hdmi2usbsoc_hdmi_out1_resetinserter_source_source_ready = hdmi2usbsoc_hdmi_out1_sink_ready;
assign hdmi2usbsoc_hdmi_out1_sink_first = hdmi2usbsoc_hdmi_out1_resetinserter_source_source_first;
assign hdmi2usbsoc_hdmi_out1_sink_last = hdmi2usbsoc_hdmi_out1_resetinserter_source_source_last;
assign hdmi2usbsoc_hdmi_out1_sink_payload_y = hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_y;
assign hdmi2usbsoc_hdmi_out1_sink_payload_cb = hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_cb;
assign hdmi2usbsoc_hdmi_out1_sink_payload_cr = hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_cr;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_valid = hdmi2usbsoc_hdmi_out1_source_valid;
assign hdmi2usbsoc_hdmi_out1_source_ready = hdmi2usbsoc_hdmi_out1_driver_sink_sink_ready;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_first = hdmi2usbsoc_hdmi_out1_source_first;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_last = hdmi2usbsoc_hdmi_out1_source_last;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_r = hdmi2usbsoc_hdmi_out1_source_payload_r;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_g = hdmi2usbsoc_hdmi_out1_source_payload_g;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_b = hdmi2usbsoc_hdmi_out1_source_payload_b;
assign hdmi2usbsoc_hdmi_out1_sink_payload_de = hdmi2usbsoc_hdmi_out1_core_source_source_param_de;
assign hdmi2usbsoc_hdmi_out1_sink_payload_vsync = hdmi2usbsoc_hdmi_out1_core_source_source_param_vsync;
assign hdmi2usbsoc_hdmi_out1_sink_payload_hsync = hdmi2usbsoc_hdmi_out1_core_source_source_param_hsync;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_de = hdmi2usbsoc_hdmi_out1_source_payload_de;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_vsync = hdmi2usbsoc_hdmi_out1_source_payload_vsync;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_hsync = hdmi2usbsoc_hdmi_out1_source_payload_hsync;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_valid = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_valid;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_sink_valid = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_valid;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_ready = hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_ready;
assign hdmi2usbsoc_hdmi_out1_core_source_source_valid = (hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_valid & ((~hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_de) | hdmi2usbsoc_hdmi_out1_core_dmareader_source_valid));

// synthesis translate_off
reg dummy_d_118;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_ready <= 1'd0;
	hdmi2usbsoc_hdmi_out1_core_dmareader_source_ready <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_out1_core_initiator_source_source_valid)) begin
		hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_ready <= 1'd1;
		hdmi2usbsoc_hdmi_out1_core_dmareader_source_ready <= 1'd1;
	end else begin
		if ((hdmi2usbsoc_hdmi_out1_core_source_source_valid & hdmi2usbsoc_hdmi_out1_core_source_source_ready)) begin
			hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_ready <= 1'd1;
			hdmi2usbsoc_hdmi_out1_core_dmareader_source_ready <= (hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_de | 1'd0);
		end
	end
// synthesis translate_off
	dummy_d_118 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hres = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hres;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hscan = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hscan;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vres = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vres;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vscan = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vscan;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_sink_payload_base = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_base;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_sink_payload_length = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_length;
assign hdmi2usbsoc_hdmi_out1_core_source_source_param_de = hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_de;
assign hdmi2usbsoc_hdmi_out1_core_source_source_param_hsync = hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_hsync;
assign hdmi2usbsoc_hdmi_out1_core_source_source_param_vsync = hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_vsync;
assign hdmi2usbsoc_hdmi_out1_core_source_source_payload_data = hdmi2usbsoc_hdmi_out1_core_dmareader_source_payload_data;
assign hdmi2usbsoc_hdmi_out1_core_i = hdmi2usbsoc_hdmi_out1_core_underflow_update_underflow_update_re;
assign hdmi2usbsoc_hdmi_out1_core_underflow_update = hdmi2usbsoc_hdmi_out1_core_o;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hres = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hscan = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vres = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vscan = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_base = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_length = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_valid = hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_valid = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_valid;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_ready = hdmi2usbsoc_hdmi_out1_core_initiator_source_source_ready;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_first = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_first;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_last = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_last;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hres = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hres;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_hscan = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hscan;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vres = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vres;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_vscan = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vscan;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_base = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_base;
assign hdmi2usbsoc_hdmi_out1_core_initiator_source_source_payload_length = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_length;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_din = {hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_last, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_first, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_length, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_base, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vscan, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vsync_end, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vsync_start, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vres, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hscan, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hsync_end, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hsync_start, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hres};
assign {hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_last, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_first, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_length, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_base, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vscan, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vsync_end, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vsync_start, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vres, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hscan, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hsync_end, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hsync_start, hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hres} = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_dout;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_ready = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_writable;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_we = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_valid;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_first = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_first;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_last = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_last;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hres = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hres;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_hscan = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_hscan;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vres = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vres;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_vscan = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_vscan;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_base = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_base;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_in_payload_length = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_sink_payload_length;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_valid = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_readable;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_first = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_first;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_last = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_last;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hres = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hres;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hsync_start;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hsync_end;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_hscan = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_hscan;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vres = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vres;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vsync_start = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vsync_start;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vsync_end = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vsync_end;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_vscan = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_vscan;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_base = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_base;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_payload_length = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_fifo_out_payload_length;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_re = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_source_ready;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_ce = (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_writable & hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_we);
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_ce = (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_readable & hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_re);
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_writable = ((hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q[1] == hdmi2usbsoc_hdmi_out1_core_initiator_cdc_consume_wdomain[1]) | (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q[0] == hdmi2usbsoc_hdmi_out1_core_initiator_cdc_consume_wdomain[0]));
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_readable = (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q != hdmi2usbsoc_hdmi_out1_core_initiator_cdc_produce_rdomain);
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_adr = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_binary[0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_dat_w = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_din;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_we = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_ce;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_rdport_adr = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary[0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_asyncfifo_dout = hdmi2usbsoc_hdmi_out1_core_initiator_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_119;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next_binary <= 2'd0;
	if (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_ce) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next_binary <= (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next_binary <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_119 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next = (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next_binary ^ hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next_binary[1]);

// synthesis translate_off
reg dummy_d_120;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary <= 2'd0;
	if (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_ce) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary <= (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_120 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next = (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary ^ hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary[1]);

// synthesis translate_off
reg dummy_d_121;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_core_timinggenerator_active <= 1'd0;
	hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_de <= 1'd0;
	hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_valid <= 1'd0;
	if (hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_valid) begin
		hdmi2usbsoc_hdmi_out1_core_timinggenerator_active <= (hdmi2usbsoc_hdmi_out1_core_timinggenerator_hactive & hdmi2usbsoc_hdmi_out1_core_timinggenerator_vactive);
		hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_valid <= 1'd1;
		if (hdmi2usbsoc_hdmi_out1_core_timinggenerator_active) begin
			hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_de <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_121 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_ready = (hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_ready & hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_last);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_base = hdmi2usbsoc_hdmi_out1_core_dmareader_sink_payload_base[31:1];
assign hdmi2usbsoc_hdmi_out1_core_dmareader_length = hdmi2usbsoc_hdmi_out1_core_dmareader_sink_payload_length[31:1];
assign hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_payload_address = (hdmi2usbsoc_hdmi_out1_core_dmareader_base + hdmi2usbsoc_hdmi_out1_core_dmareader_offset);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_valid = hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_valid;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_ready = hdmi2usbsoc_hdmi_out1_core_dmareader_source_ready;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_first = hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_first;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_last = hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_last;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_payload_data = hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_payload_data;
assign hdmi2usbsoc_litedramport3_cmd_payload_we1 = 1'd0;
assign hdmi2usbsoc_litedramport3_cmd_valid1 = (hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_valid & hdmi2usbsoc_hdmi_out1_core_dmareader_request_enable);
assign hdmi2usbsoc_litedramport3_cmd_payload_adr1 = hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_payload_address;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_ready = (hdmi2usbsoc_litedramport3_cmd_ready1 & hdmi2usbsoc_hdmi_out1_core_dmareader_request_enable);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_request_issued = (hdmi2usbsoc_litedramport3_cmd_valid1 & hdmi2usbsoc_litedramport3_cmd_ready1);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_request_enable = (hdmi2usbsoc_hdmi_out1_core_dmareader_rsv_level != 13'd4096);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_valid = hdmi2usbsoc_litedramport3_rdata_valid1;
assign hdmi2usbsoc_litedramport3_rdata_ready1 = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_ready;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_first = hdmi2usbsoc_litedramport3_rdata_first1;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_last = hdmi2usbsoc_litedramport3_rdata_last1;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_payload_data = hdmi2usbsoc_litedramport3_rdata_payload_data1;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_valid = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_valid;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_ready = hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_ready;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_first = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_first;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_last = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_last;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_payload_data = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_data_dequeued = (hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_valid & hdmi2usbsoc_hdmi_out1_core_dmareader_source_source_ready);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_ready = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_valid = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_readable;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_first = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_last = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_payload_data = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_re = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_source_ready;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_re = (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_readable & ((~hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_readable) | hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_re));
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level1 = (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 + hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_readable);

// synthesis translate_off
reg dummy_d_122;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_adr <= 12'd0;
	if (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_replace) begin
		hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_produce;
	end
// synthesis translate_off
	dummy_d_122 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_we = (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_replace));
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_do_read = (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_adr = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_consume;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_re = hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_do_read;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 != 13'd4096);
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 != 1'd0);

// synthesis translate_off
reg dummy_d_123;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_valid <= 1'd0;
	videoout1_next_state <= 1'd0;
	hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value <= 26'd0;
	hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value_ce <= 1'd0;
	hdmi2usbsoc_hdmi_out1_core_dmareader_sink_ready <= 1'd0;
	hdmi2usbsoc_litedramport3_flush <= 1'd0;
	videoout1_next_state <= videoout1_state;
	case (videoout1_state)
		1'd1: begin
			hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_valid <= 1'd1;
			if (hdmi2usbsoc_hdmi_out1_core_dmareader_sink_sink_ready) begin
				hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value <= (hdmi2usbsoc_hdmi_out1_core_dmareader_offset + 1'd1);
				hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value_ce <= 1'd1;
				if ((hdmi2usbsoc_hdmi_out1_core_dmareader_offset == (hdmi2usbsoc_hdmi_out1_core_dmareader_length - 1'd1))) begin
					hdmi2usbsoc_hdmi_out1_core_dmareader_sink_ready <= 1'd1;
					videoout1_next_state <= 1'd0;
				end
			end
		end
		default: begin
			hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value <= 1'd0;
			hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value_ce <= 1'd1;
			if (hdmi2usbsoc_hdmi_out1_core_dmareader_sink_valid) begin
				videoout1_next_state <= 1'd1;
			end else begin
				hdmi2usbsoc_litedramport3_flush <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_123 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_core_o = (hdmi2usbsoc_hdmi_out1_core_toggle_o ^ hdmi2usbsoc_hdmi_out1_core_toggle_o_r);
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe = hdmi2usbsoc_hdmi_out1_driver_clocking_serdesstrobe;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_valid = hdmi2usbsoc_hdmi_out1_driver_sink_sink_valid;
assign hdmi2usbsoc_hdmi_out1_driver_sink_sink_ready = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_ready;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_first = hdmi2usbsoc_hdmi_out1_driver_sink_sink_first;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_last = hdmi2usbsoc_hdmi_out1_driver_sink_sink_last;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_r = hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_r;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_g = hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_g;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_b = hdmi2usbsoc_hdmi_out1_driver_sink_sink_payload_b;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_hsync = hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_hsync;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_vsync = hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_vsync;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_de = hdmi2usbsoc_hdmi_out1_driver_sink_sink_param_de;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_ready = 1'd1;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0 = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_b;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0 = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_g;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0 = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_payload_r;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_c = {hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_vsync, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_hsync};
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_c = 1'd0;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_c = 1'd0;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_de = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_de;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_de = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_de;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_de = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_sink_param_de;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x_pol;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n = ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1d > 3'd4) | ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1d == 3'd4) & (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0])));
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x_pol;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n = ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1d > 3'd4) | ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1d == 3'd4) & (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0])));
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x = hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x_pol;
assign hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n = ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1d > 3'd4) | ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1d == 3'd4) & (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0])));

// synthesis translate_off
reg dummy_d_124;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready <= 1'd0;
	hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_payload_data <= 8'd0;
	hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_payload_data <= 8'd0;
	hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_payload_data <= 8'd0;
	hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_valid <= 1'd0;
	hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_valid <= 1'd0;
	hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_valid <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_out1_resetinserter_parity_in)) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_y;
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_cb_cr;
		hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready <= (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_ready & hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_ready);
	end else begin
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_y;
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_valid <= (hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready);
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_payload_data <= hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_payload_cb_cr;
		hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready <= (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_ready & hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_ready);
	end
// synthesis translate_off
	dummy_d_124 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_resetinserter_source_source_valid = ((hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_valid & hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_valid) & hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_valid);
assign hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_y = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_cb = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_source_source_payload_cr = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_ready = (hdmi2usbsoc_hdmi_out1_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out1_resetinserter_source_source_ready);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_ready = ((hdmi2usbsoc_hdmi_out1_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out1_resetinserter_source_source_ready) & hdmi2usbsoc_hdmi_out1_resetinserter_parity_out);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_ready = ((hdmi2usbsoc_hdmi_out1_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out1_resetinserter_source_source_ready) & hdmi2usbsoc_hdmi_out1_resetinserter_parity_out);
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_ready = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_valid = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_first = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_last = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_payload_data = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_re = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_source_ready;

// synthesis translate_off
reg dummy_d_125;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_replace) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_produce;
	end
// synthesis translate_off
	dummy_d_125 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_we = (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_replace));
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_do_read = (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_rdport_adr = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_consume;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level != 3'd4);
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_ready = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_valid = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_first = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_last = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_payload_data = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_re = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_source_ready;

// synthesis translate_off
reg dummy_d_126;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_replace) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_produce;
	end
// synthesis translate_off
	dummy_d_126 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_we = (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_replace));
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_do_read = (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_rdport_adr = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_consume;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level != 3'd4);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_din = {hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_last, hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_first, hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_payload_data};
assign {hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_last, hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_first, hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_payload_data} = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_dout;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_ready = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_writable;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_we = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_valid;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_first = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_first;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_last = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_last;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_in_payload_data = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_sink_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_valid = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_readable;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_first = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_first;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_last = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_last;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_payload_data = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_fifo_out_payload_data;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_re = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_source_ready;

// synthesis translate_off
reg dummy_d_127;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_adr <= 2'd0;
	if (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_replace) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_adr <= (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_produce - 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_adr <= hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_produce;
	end
// synthesis translate_off
	dummy_d_127 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_dat_w = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_din;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_we = (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_we & (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_writable | hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_replace));
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_do_read = (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_readable & hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_re);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_rdport_adr = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_consume;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_dout = hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_rdport_dat_r;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_writable = (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level != 3'd4);
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_readable = (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level != 1'd0);
assign hdmi2usbsoc_hdmi_out1_pipe_ce = (hdmi2usbsoc_hdmi_out1_source_ready | (~hdmi2usbsoc_hdmi_out1_valid_n3));
assign hdmi2usbsoc_hdmi_out1_sink_ready = hdmi2usbsoc_hdmi_out1_pipe_ce;
assign hdmi2usbsoc_hdmi_out1_source_valid = hdmi2usbsoc_hdmi_out1_valid_n3;
assign hdmi2usbsoc_hdmi_out1_busy = ((((1'd0 | hdmi2usbsoc_hdmi_out1_valid_n0) | hdmi2usbsoc_hdmi_out1_valid_n1) | hdmi2usbsoc_hdmi_out1_valid_n2) | hdmi2usbsoc_hdmi_out1_valid_n3);
assign hdmi2usbsoc_hdmi_out1_source_first = hdmi2usbsoc_hdmi_out1_first_n3;
assign hdmi2usbsoc_hdmi_out1_source_last = hdmi2usbsoc_hdmi_out1_last_n3;
assign hdmi2usbsoc_hdmi_out1_ce = hdmi2usbsoc_hdmi_out1_pipe_ce;
assign hdmi2usbsoc_hdmi_out1_sink_y = hdmi2usbsoc_hdmi_out1_sink_payload_y;
assign hdmi2usbsoc_hdmi_out1_sink_cb = hdmi2usbsoc_hdmi_out1_sink_payload_cb;
assign hdmi2usbsoc_hdmi_out1_sink_cr = hdmi2usbsoc_hdmi_out1_sink_payload_cr;
assign hdmi2usbsoc_hdmi_out1_source_payload_r = hdmi2usbsoc_hdmi_out1_source_r;
assign hdmi2usbsoc_hdmi_out1_source_payload_g = hdmi2usbsoc_hdmi_out1_source_g;
assign hdmi2usbsoc_hdmi_out1_source_payload_b = hdmi2usbsoc_hdmi_out1_source_b;
assign hdmi2usbsoc_hdmi_out1_source_payload_hsync = hdmi2usbsoc_hdmi_out1_next_s5;
assign hdmi2usbsoc_hdmi_out1_source_payload_vsync = hdmi2usbsoc_hdmi_out1_next_s11;
assign hdmi2usbsoc_hdmi_out1_source_payload_de = hdmi2usbsoc_hdmi_out1_next_s17;
assign encoder_reader_source_valid = encoder_reader_source_source_valid;
assign encoder_reader_source_source_ready = encoder_reader_source_ready;
assign encoder_reader_source_first = encoder_reader_source_source_first;
assign encoder_reader_source_last = encoder_reader_source_source_last;
assign encoder_reader_source_payload_data = encoder_reader_source_source_payload_data;
assign encoder_reader_h_next = (encoder_reader_h + 4'd8);
assign encoder_reader_read_address = ((encoder_reader_v * encoder_reader_h_width_storage) + encoder_reader_h);
assign encoder_reader_sink_sink_payload_address = (encoder_reader_base[31:4] + encoder_reader_read_address[26:3]);
assign encoder_port_new_port_cmd_payload_we = 1'd0;
assign encoder_port_new_port_cmd_valid = (encoder_reader_sink_sink_valid & encoder_reader_request_enable);
assign encoder_port_new_port_cmd_payload_adr = encoder_reader_sink_sink_payload_address;
assign encoder_reader_sink_sink_ready = (encoder_port_new_port_cmd_ready & encoder_reader_request_enable);
assign encoder_reader_request_issued = (encoder_port_new_port_cmd_valid & encoder_port_new_port_cmd_ready);
assign encoder_reader_request_enable = (encoder_reader_rsv_level != 5'd16);
assign encoder_reader_fifo_sink_valid = encoder_port_new_port_rdata_valid;
assign encoder_port_new_port_rdata_ready = encoder_reader_fifo_sink_ready;
assign encoder_reader_fifo_sink_first = encoder_port_new_port_rdata_first;
assign encoder_reader_fifo_sink_last = encoder_port_new_port_rdata_last;
assign encoder_reader_fifo_sink_payload_data = encoder_port_new_port_rdata_payload_data;
assign encoder_reader_source_source_valid = encoder_reader_fifo_source_valid;
assign encoder_reader_fifo_source_ready = encoder_reader_source_source_ready;
assign encoder_reader_source_source_first = encoder_reader_fifo_source_first;
assign encoder_reader_source_source_last = encoder_reader_fifo_source_last;
assign encoder_reader_source_source_payload_data = encoder_reader_fifo_source_payload_data;
assign encoder_reader_data_dequeued = (encoder_reader_source_source_valid & encoder_reader_source_source_ready);
assign encoder_reader_fifo_syncfifo_din = {encoder_reader_fifo_fifo_in_last, encoder_reader_fifo_fifo_in_first, encoder_reader_fifo_fifo_in_payload_data};
assign {encoder_reader_fifo_fifo_out_last, encoder_reader_fifo_fifo_out_first, encoder_reader_fifo_fifo_out_payload_data} = encoder_reader_fifo_syncfifo_dout;
assign encoder_reader_fifo_sink_ready = encoder_reader_fifo_syncfifo_writable;
assign encoder_reader_fifo_syncfifo_we = encoder_reader_fifo_sink_valid;
assign encoder_reader_fifo_fifo_in_first = encoder_reader_fifo_sink_first;
assign encoder_reader_fifo_fifo_in_last = encoder_reader_fifo_sink_last;
assign encoder_reader_fifo_fifo_in_payload_data = encoder_reader_fifo_sink_payload_data;
assign encoder_reader_fifo_source_valid = encoder_reader_fifo_syncfifo_readable;
assign encoder_reader_fifo_source_first = encoder_reader_fifo_fifo_out_first;
assign encoder_reader_fifo_source_last = encoder_reader_fifo_fifo_out_last;
assign encoder_reader_fifo_source_payload_data = encoder_reader_fifo_fifo_out_payload_data;
assign encoder_reader_fifo_syncfifo_re = encoder_reader_fifo_source_ready;

// synthesis translate_off
reg dummy_d_128;
// synthesis translate_on
always @(*) begin
	encoder_reader_fifo_wrport_adr <= 4'd0;
	if (encoder_reader_fifo_replace) begin
		encoder_reader_fifo_wrport_adr <= (encoder_reader_fifo_produce - 1'd1);
	end else begin
		encoder_reader_fifo_wrport_adr <= encoder_reader_fifo_produce;
	end
// synthesis translate_off
	dummy_d_128 <= dummy_s;
// synthesis translate_on
end
assign encoder_reader_fifo_wrport_dat_w = encoder_reader_fifo_syncfifo_din;
assign encoder_reader_fifo_wrport_we = (encoder_reader_fifo_syncfifo_we & (encoder_reader_fifo_syncfifo_writable | encoder_reader_fifo_replace));
assign encoder_reader_fifo_do_read = (encoder_reader_fifo_syncfifo_readable & encoder_reader_fifo_syncfifo_re);
assign encoder_reader_fifo_rdport_adr = encoder_reader_fifo_consume;
assign encoder_reader_fifo_syncfifo_dout = encoder_reader_fifo_rdport_dat_r;
assign encoder_reader_fifo_syncfifo_writable = (encoder_reader_fifo_level != 5'd16);
assign encoder_reader_fifo_syncfifo_readable = (encoder_reader_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_129;
// synthesis translate_on
always @(*) begin
	encoderdmareader_next_state <= 1'd0;
	encoder_reader_status <= 1'd0;
	encoder_reader_sink_sink_valid <= 1'd0;
	encoder_reader_h_clr <= 1'd0;
	encoder_reader_h_clr_lsb <= 1'd0;
	encoder_reader_h_inc <= 1'd0;
	encoder_reader_v_clr <= 1'd0;
	encoder_reader_v_inc <= 1'd0;
	encoder_reader_v_dec7 <= 1'd0;
	encoderdmareader_next_state <= encoderdmareader_state;
	case (encoderdmareader_state)
		1'd1: begin
			encoder_reader_sink_sink_valid <= 1'd1;
			if (encoder_reader_sink_sink_ready) begin
				if ((encoder_reader_h_next[2:0] == 1'd0)) begin
					if ((encoder_reader_v[2:0] == 3'd7)) begin
						if ((encoder_reader_h >= (encoder_reader_h_width_storage - 4'd8))) begin
							encoder_reader_h_clr <= 1'd1;
							encoder_reader_v_inc <= 1'd1;
							if ((encoder_reader_v >= (encoder_reader_v_width_storage - 1'd1))) begin
								encoderdmareader_next_state <= 1'd0;
							end
						end else begin
							encoder_reader_h_inc <= 1'd1;
							encoder_reader_v_dec7 <= 1'd1;
						end
					end else begin
						encoder_reader_h_clr_lsb <= 1'd1;
						encoder_reader_v_inc <= 1'd1;
					end
				end else begin
					encoder_reader_h_inc <= 1'd1;
				end
			end
		end
		default: begin
			encoder_reader_h_clr <= 1'd1;
			encoder_reader_v_clr <= 1'd1;
			if ((encoder_reader_start_r & encoder_reader_start_re)) begin
				encoderdmareader_next_state <= 1'd1;
			end else begin
				encoder_reader_status <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_129 <= dummy_s;
// synthesis translate_on
end
assign encoder_cdc_asyncfifo_din = {encoder_cdc_fifo_in_last, encoder_cdc_fifo_in_first, encoder_cdc_fifo_in_payload_data};
assign {encoder_cdc_fifo_out_last, encoder_cdc_fifo_out_first, encoder_cdc_fifo_out_payload_data} = encoder_cdc_asyncfifo_dout;
assign encoder_cdc_sink_ready = encoder_cdc_asyncfifo_writable;
assign encoder_cdc_asyncfifo_we = encoder_cdc_sink_valid;
assign encoder_cdc_fifo_in_first = encoder_cdc_sink_first;
assign encoder_cdc_fifo_in_last = encoder_cdc_sink_last;
assign encoder_cdc_fifo_in_payload_data = encoder_cdc_sink_payload_data;
assign encoder_cdc_source_valid = encoder_cdc_asyncfifo_readable;
assign encoder_cdc_source_first = encoder_cdc_fifo_out_first;
assign encoder_cdc_source_last = encoder_cdc_fifo_out_last;
assign encoder_cdc_source_payload_data = encoder_cdc_fifo_out_payload_data;
assign encoder_cdc_asyncfifo_re = encoder_cdc_source_ready;
assign encoder_cdc_graycounter0_ce = (encoder_cdc_asyncfifo_writable & encoder_cdc_asyncfifo_we);
assign encoder_cdc_graycounter1_ce = (encoder_cdc_asyncfifo_readable & encoder_cdc_asyncfifo_re);
assign encoder_cdc_asyncfifo_writable = (((encoder_cdc_graycounter0_q[2] == encoder_cdc_consume_wdomain[2]) | (encoder_cdc_graycounter0_q[1] == encoder_cdc_consume_wdomain[1])) | (encoder_cdc_graycounter0_q[0] != encoder_cdc_consume_wdomain[0]));
assign encoder_cdc_asyncfifo_readable = (encoder_cdc_graycounter1_q != encoder_cdc_produce_rdomain);
assign encoder_cdc_wrport_adr = encoder_cdc_graycounter0_q_binary[1:0];
assign encoder_cdc_wrport_dat_w = encoder_cdc_asyncfifo_din;
assign encoder_cdc_wrport_we = encoder_cdc_graycounter0_ce;
assign encoder_cdc_rdport_adr = encoder_cdc_graycounter1_q_next_binary[1:0];
assign encoder_cdc_asyncfifo_dout = encoder_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_130;
// synthesis translate_on
always @(*) begin
	encoder_cdc_graycounter0_q_next_binary <= 3'd0;
	if (encoder_cdc_graycounter0_ce) begin
		encoder_cdc_graycounter0_q_next_binary <= (encoder_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		encoder_cdc_graycounter0_q_next_binary <= encoder_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_130 <= dummy_s;
// synthesis translate_on
end
assign encoder_cdc_graycounter0_q_next = (encoder_cdc_graycounter0_q_next_binary ^ encoder_cdc_graycounter0_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_131;
// synthesis translate_on
always @(*) begin
	encoder_cdc_graycounter1_q_next_binary <= 3'd0;
	if (encoder_cdc_graycounter1_ce) begin
		encoder_cdc_graycounter1_q_next_binary <= (encoder_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		encoder_cdc_graycounter1_q_next_binary <= encoder_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_131 <= dummy_s;
// synthesis translate_on
end
assign encoder_cdc_graycounter1_q_next = (encoder_cdc_graycounter1_q_next_binary ^ encoder_cdc_graycounter1_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_132;
// synthesis translate_on
always @(*) begin
	encoderbuffer_write_port_adr <= 4'd0;
	encoderbuffer_write_port_adr <= encoderbuffer_v_write;
	encoderbuffer_write_port_adr[3] <= encoderbuffer_write_sel;
// synthesis translate_off
	dummy_d_132 <= dummy_s;
// synthesis translate_on
end
assign encoderbuffer_write_port_dat_w = encoderbuffer_sink_payload_data;
assign encoderbuffer_write_port_we = (encoderbuffer_sink_valid & encoderbuffer_sink_ready);

// synthesis translate_off
reg dummy_d_133;
// synthesis translate_on
always @(*) begin
	encoderbuffer_read_port_adr <= 4'd0;
	encoderbuffer_read_port_adr <= encoderbuffer_v_read;
	encoderbuffer_read_port_adr[3] <= encoderbuffer_read_sel;
// synthesis translate_off
	dummy_d_133 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_134;
// synthesis translate_on
always @(*) begin
	encoderbuffer_source_payload_data <= 16'd0;
	case (encoderbuffer_h_read)
		1'd0: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[127:112];
		end
		1'd1: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[111:96];
		end
		2'd2: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[95:80];
		end
		2'd3: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[79:64];
		end
		3'd4: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[63:48];
		end
		3'd5: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[47:32];
		end
		3'd6: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[31:16];
		end
		default: begin
			encoderbuffer_source_payload_data <= encoderbuffer_read_port_dat_r[15:0];
		end
	endcase
// synthesis translate_off
	dummy_d_134 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_135;
// synthesis translate_on
always @(*) begin
	encoderbuffer_sink_ready <= 1'd0;
	encoderbuffer_write_swap <= 1'd0;
	encoderbuffer_v_write_clr <= 1'd0;
	encoderbuffer_v_write_inc <= 1'd0;
	fsm0_next_state <= 1'd0;
	fsm0_next_state <= fsm0_state;
	case (fsm0_state)
		1'd1: begin
			encoderbuffer_sink_ready <= 1'd1;
			if (encoderbuffer_sink_valid) begin
				if ((encoderbuffer_v_write == 3'd7)) begin
					encoderbuffer_write_swap <= 1'd1;
					fsm0_next_state <= 1'd0;
				end else begin
					encoderbuffer_v_write_inc <= 1'd1;
				end
			end
		end
		default: begin
			encoderbuffer_v_write_clr <= 1'd1;
			if ((encoderbuffer_write_sel != encoderbuffer_read_sel)) begin
				fsm0_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_135 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_136;
// synthesis translate_on
always @(*) begin
	encoderbuffer_h_read_clr <= 1'd0;
	encoderbuffer_h_read_inc <= 1'd0;
	encoderbuffer_source_valid <= 1'd0;
	encoderbuffer_v_read_clr <= 1'd0;
	encoderbuffer_v_read_inc <= 1'd0;
	encoderbuffer_source_last <= 1'd0;
	fsm1_next_state <= 1'd0;
	encoderbuffer_read_swap <= 1'd0;
	fsm1_next_state <= fsm1_state;
	case (fsm1_state)
		1'd1: begin
			encoderbuffer_source_valid <= 1'd1;
			encoderbuffer_source_last <= ((encoderbuffer_h_read == 3'd7) & (encoderbuffer_v_read == 3'd7));
			if (encoderbuffer_source_ready) begin
				if ((encoderbuffer_h_read == 3'd7)) begin
					encoderbuffer_h_read_clr <= 1'd1;
					if ((encoderbuffer_v_read == 3'd7)) begin
						fsm1_next_state <= 1'd0;
					end else begin
						encoderbuffer_v_read_inc <= 1'd1;
					end
				end else begin
					encoderbuffer_h_read_inc <= 1'd1;
				end
			end
		end
		default: begin
			encoderbuffer_h_read_clr <= 1'd1;
			encoderbuffer_v_read_clr <= 1'd1;
			if ((encoderbuffer_read_sel == encoderbuffer_write_sel)) begin
				encoderbuffer_read_swap <= 1'd1;
				fsm1_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_136 <= dummy_s;
// synthesis translate_on
end
assign encoder_sink_sink_valid1 = encoder_sink_sink_valid0;
assign encoder_sink_sink_ready0 = encoder_sink_sink_ready1;
assign encoder_sink_sink_first1 = encoder_sink_sink_first0;
assign encoder_sink_sink_last1 = encoder_sink_sink_last0;
assign encoder_sink_sink_payload_y = encoder_sink_sink_payload_data[7:0];
assign encoder_sink_sink_payload_cb_cr = encoder_sink_sink_payload_data[15:8];
assign encoder_fdct_fifo_q = encoder_fdct_data_d4;
assign encoder_fdct_fifo_hf_full = encoder_source_source_valid1;
assign encoder_source_source_ready1 = encoder_fdct_fifo_rd;
assign encoder_output_fifo_almost_full = (encoder_output_fifo_level1 > 10'd896);
assign encoder_source_source_valid0 = encoder_output_fifo_source_valid;
assign encoder_output_fifo_source_ready = encoder_source_source_ready0;
assign encoder_source_source_first = encoder_output_fifo_source_first;
assign encoder_source_source_last = encoder_output_fifo_source_last;
assign encoder_source_source_payload_data = encoder_output_fifo_source_payload_data;

// synthesis translate_off
reg dummy_d_137;
// synthesis translate_on
always @(*) begin
	encoder_y_fifo_sink_payload_data <= 8'd0;
	encoder_cb_fifo_sink_payload_data <= 8'd0;
	encoder_sink_sink_ready1 <= 1'd0;
	encoder_cr_fifo_sink_payload_data <= 8'd0;
	encoder_y_fifo_sink_valid <= 1'd0;
	encoder_cb_fifo_sink_valid <= 1'd0;
	encoder_cr_fifo_sink_valid <= 1'd0;
	if ((~encoder_parity_in)) begin
		encoder_y_fifo_sink_valid <= (encoder_sink_sink_valid1 & encoder_sink_sink_ready1);
		encoder_y_fifo_sink_payload_data <= encoder_sink_sink_payload_y;
		encoder_cb_fifo_sink_valid <= (encoder_sink_sink_valid1 & encoder_sink_sink_ready1);
		encoder_cb_fifo_sink_payload_data <= encoder_sink_sink_payload_cb_cr;
		encoder_sink_sink_ready1 <= (encoder_y_fifo_sink_ready & encoder_cb_fifo_sink_ready);
	end else begin
		encoder_y_fifo_sink_valid <= (encoder_sink_sink_valid1 & encoder_sink_sink_ready1);
		encoder_y_fifo_sink_payload_data <= encoder_sink_sink_payload_y;
		encoder_cr_fifo_sink_valid <= (encoder_sink_sink_valid1 & encoder_sink_sink_ready1);
		encoder_cr_fifo_sink_payload_data <= encoder_sink_sink_payload_cb_cr;
		encoder_sink_sink_ready1 <= (encoder_y_fifo_sink_ready & encoder_cr_fifo_sink_ready);
	end
// synthesis translate_off
	dummy_d_137 <= dummy_s;
// synthesis translate_on
end
assign encoder_source_source_valid1 = ((encoder_y_fifo_source_valid & encoder_cb_fifo_source_valid) & encoder_cr_fifo_source_valid);
assign encoder_source_source_payload_y = encoder_y_fifo_source_payload_data;
assign encoder_source_source_payload_cb = encoder_cb_fifo_source_payload_data;
assign encoder_source_source_payload_cr = encoder_cr_fifo_source_payload_data;
assign encoder_y_fifo_source_ready = (encoder_source_source_valid1 & encoder_source_source_ready1);
assign encoder_cb_fifo_source_ready = ((encoder_source_source_valid1 & encoder_source_source_ready1) & encoder_parity_out);
assign encoder_cr_fifo_source_ready = ((encoder_source_source_valid1 & encoder_source_source_ready1) & encoder_parity_out);
assign encoder_y_fifo_syncfifo_din = {encoder_y_fifo_fifo_in_last, encoder_y_fifo_fifo_in_first, encoder_y_fifo_fifo_in_payload_data};
assign {encoder_y_fifo_fifo_out_last, encoder_y_fifo_fifo_out_first, encoder_y_fifo_fifo_out_payload_data} = encoder_y_fifo_syncfifo_dout;
assign encoder_y_fifo_sink_ready = encoder_y_fifo_syncfifo_writable;
assign encoder_y_fifo_syncfifo_we = encoder_y_fifo_sink_valid;
assign encoder_y_fifo_fifo_in_first = encoder_y_fifo_sink_first;
assign encoder_y_fifo_fifo_in_last = encoder_y_fifo_sink_last;
assign encoder_y_fifo_fifo_in_payload_data = encoder_y_fifo_sink_payload_data;
assign encoder_y_fifo_source_valid = encoder_y_fifo_syncfifo_readable;
assign encoder_y_fifo_source_first = encoder_y_fifo_fifo_out_first;
assign encoder_y_fifo_source_last = encoder_y_fifo_fifo_out_last;
assign encoder_y_fifo_source_payload_data = encoder_y_fifo_fifo_out_payload_data;
assign encoder_y_fifo_syncfifo_re = encoder_y_fifo_source_ready;

// synthesis translate_off
reg dummy_d_138;
// synthesis translate_on
always @(*) begin
	encoder_y_fifo_wrport_adr <= 2'd0;
	if (encoder_y_fifo_replace) begin
		encoder_y_fifo_wrport_adr <= (encoder_y_fifo_produce - 1'd1);
	end else begin
		encoder_y_fifo_wrport_adr <= encoder_y_fifo_produce;
	end
// synthesis translate_off
	dummy_d_138 <= dummy_s;
// synthesis translate_on
end
assign encoder_y_fifo_wrport_dat_w = encoder_y_fifo_syncfifo_din;
assign encoder_y_fifo_wrport_we = (encoder_y_fifo_syncfifo_we & (encoder_y_fifo_syncfifo_writable | encoder_y_fifo_replace));
assign encoder_y_fifo_do_read = (encoder_y_fifo_syncfifo_readable & encoder_y_fifo_syncfifo_re);
assign encoder_y_fifo_rdport_adr = encoder_y_fifo_consume;
assign encoder_y_fifo_syncfifo_dout = encoder_y_fifo_rdport_dat_r;
assign encoder_y_fifo_syncfifo_writable = (encoder_y_fifo_level != 3'd4);
assign encoder_y_fifo_syncfifo_readable = (encoder_y_fifo_level != 1'd0);
assign encoder_cb_fifo_syncfifo_din = {encoder_cb_fifo_fifo_in_last, encoder_cb_fifo_fifo_in_first, encoder_cb_fifo_fifo_in_payload_data};
assign {encoder_cb_fifo_fifo_out_last, encoder_cb_fifo_fifo_out_first, encoder_cb_fifo_fifo_out_payload_data} = encoder_cb_fifo_syncfifo_dout;
assign encoder_cb_fifo_sink_ready = encoder_cb_fifo_syncfifo_writable;
assign encoder_cb_fifo_syncfifo_we = encoder_cb_fifo_sink_valid;
assign encoder_cb_fifo_fifo_in_first = encoder_cb_fifo_sink_first;
assign encoder_cb_fifo_fifo_in_last = encoder_cb_fifo_sink_last;
assign encoder_cb_fifo_fifo_in_payload_data = encoder_cb_fifo_sink_payload_data;
assign encoder_cb_fifo_source_valid = encoder_cb_fifo_syncfifo_readable;
assign encoder_cb_fifo_source_first = encoder_cb_fifo_fifo_out_first;
assign encoder_cb_fifo_source_last = encoder_cb_fifo_fifo_out_last;
assign encoder_cb_fifo_source_payload_data = encoder_cb_fifo_fifo_out_payload_data;
assign encoder_cb_fifo_syncfifo_re = encoder_cb_fifo_source_ready;

// synthesis translate_off
reg dummy_d_139;
// synthesis translate_on
always @(*) begin
	encoder_cb_fifo_wrport_adr <= 2'd0;
	if (encoder_cb_fifo_replace) begin
		encoder_cb_fifo_wrport_adr <= (encoder_cb_fifo_produce - 1'd1);
	end else begin
		encoder_cb_fifo_wrport_adr <= encoder_cb_fifo_produce;
	end
// synthesis translate_off
	dummy_d_139 <= dummy_s;
// synthesis translate_on
end
assign encoder_cb_fifo_wrport_dat_w = encoder_cb_fifo_syncfifo_din;
assign encoder_cb_fifo_wrport_we = (encoder_cb_fifo_syncfifo_we & (encoder_cb_fifo_syncfifo_writable | encoder_cb_fifo_replace));
assign encoder_cb_fifo_do_read = (encoder_cb_fifo_syncfifo_readable & encoder_cb_fifo_syncfifo_re);
assign encoder_cb_fifo_rdport_adr = encoder_cb_fifo_consume;
assign encoder_cb_fifo_syncfifo_dout = encoder_cb_fifo_rdport_dat_r;
assign encoder_cb_fifo_syncfifo_writable = (encoder_cb_fifo_level != 3'd4);
assign encoder_cb_fifo_syncfifo_readable = (encoder_cb_fifo_level != 1'd0);
assign encoder_cr_fifo_syncfifo_din = {encoder_cr_fifo_fifo_in_last, encoder_cr_fifo_fifo_in_first, encoder_cr_fifo_fifo_in_payload_data};
assign {encoder_cr_fifo_fifo_out_last, encoder_cr_fifo_fifo_out_first, encoder_cr_fifo_fifo_out_payload_data} = encoder_cr_fifo_syncfifo_dout;
assign encoder_cr_fifo_sink_ready = encoder_cr_fifo_syncfifo_writable;
assign encoder_cr_fifo_syncfifo_we = encoder_cr_fifo_sink_valid;
assign encoder_cr_fifo_fifo_in_first = encoder_cr_fifo_sink_first;
assign encoder_cr_fifo_fifo_in_last = encoder_cr_fifo_sink_last;
assign encoder_cr_fifo_fifo_in_payload_data = encoder_cr_fifo_sink_payload_data;
assign encoder_cr_fifo_source_valid = encoder_cr_fifo_syncfifo_readable;
assign encoder_cr_fifo_source_first = encoder_cr_fifo_fifo_out_first;
assign encoder_cr_fifo_source_last = encoder_cr_fifo_fifo_out_last;
assign encoder_cr_fifo_source_payload_data = encoder_cr_fifo_fifo_out_payload_data;
assign encoder_cr_fifo_syncfifo_re = encoder_cr_fifo_source_ready;

// synthesis translate_off
reg dummy_d_140;
// synthesis translate_on
always @(*) begin
	encoder_cr_fifo_wrport_adr <= 2'd0;
	if (encoder_cr_fifo_replace) begin
		encoder_cr_fifo_wrport_adr <= (encoder_cr_fifo_produce - 1'd1);
	end else begin
		encoder_cr_fifo_wrport_adr <= encoder_cr_fifo_produce;
	end
// synthesis translate_off
	dummy_d_140 <= dummy_s;
// synthesis translate_on
end
assign encoder_cr_fifo_wrport_dat_w = encoder_cr_fifo_syncfifo_din;
assign encoder_cr_fifo_wrport_we = (encoder_cr_fifo_syncfifo_we & (encoder_cr_fifo_syncfifo_writable | encoder_cr_fifo_replace));
assign encoder_cr_fifo_do_read = (encoder_cr_fifo_syncfifo_readable & encoder_cr_fifo_syncfifo_re);
assign encoder_cr_fifo_rdport_adr = encoder_cr_fifo_consume;
assign encoder_cr_fifo_syncfifo_dout = encoder_cr_fifo_rdport_dat_r;
assign encoder_cr_fifo_syncfifo_writable = (encoder_cr_fifo_level != 3'd4);
assign encoder_cr_fifo_syncfifo_readable = (encoder_cr_fifo_level != 1'd0);
assign encoder_output_fifo_syncfifo_din = {encoder_output_fifo_fifo_in_last, encoder_output_fifo_fifo_in_first, encoder_output_fifo_fifo_in_payload_data};
assign {encoder_output_fifo_fifo_out_last, encoder_output_fifo_fifo_out_first, encoder_output_fifo_fifo_out_payload_data} = encoder_output_fifo_syncfifo_dout;
assign encoder_output_fifo_sink_ready = encoder_output_fifo_syncfifo_writable;
assign encoder_output_fifo_syncfifo_we = encoder_output_fifo_sink_valid;
assign encoder_output_fifo_fifo_in_first = encoder_output_fifo_sink_first;
assign encoder_output_fifo_fifo_in_last = encoder_output_fifo_sink_last;
assign encoder_output_fifo_fifo_in_payload_data = encoder_output_fifo_sink_payload_data;
assign encoder_output_fifo_source_valid = encoder_output_fifo_readable;
assign encoder_output_fifo_source_first = encoder_output_fifo_fifo_out_first;
assign encoder_output_fifo_source_last = encoder_output_fifo_fifo_out_last;
assign encoder_output_fifo_source_payload_data = encoder_output_fifo_fifo_out_payload_data;
assign encoder_output_fifo_re = encoder_output_fifo_source_ready;
assign encoder_output_fifo_syncfifo_re = (encoder_output_fifo_syncfifo_readable & ((~encoder_output_fifo_readable) | encoder_output_fifo_re));
assign encoder_output_fifo_level1 = (encoder_output_fifo_level0 + encoder_output_fifo_readable);

// synthesis translate_off
reg dummy_d_141;
// synthesis translate_on
always @(*) begin
	encoder_output_fifo_wrport_adr <= 10'd0;
	if (encoder_output_fifo_replace) begin
		encoder_output_fifo_wrport_adr <= (encoder_output_fifo_produce - 1'd1);
	end else begin
		encoder_output_fifo_wrport_adr <= encoder_output_fifo_produce;
	end
// synthesis translate_off
	dummy_d_141 <= dummy_s;
// synthesis translate_on
end
assign encoder_output_fifo_wrport_dat_w = encoder_output_fifo_syncfifo_din;
assign encoder_output_fifo_wrport_we = (encoder_output_fifo_syncfifo_we & (encoder_output_fifo_syncfifo_writable | encoder_output_fifo_replace));
assign encoder_output_fifo_do_read = (encoder_output_fifo_syncfifo_readable & encoder_output_fifo_syncfifo_re);
assign encoder_output_fifo_rdport_adr = encoder_output_fifo_consume;
assign encoder_output_fifo_syncfifo_dout = encoder_output_fifo_rdport_dat_r;
assign encoder_output_fifo_rdport_re = encoder_output_fifo_do_read;
assign encoder_output_fifo_syncfifo_writable = (encoder_output_fifo_level0 != 11'd1024);
assign encoder_output_fifo_syncfifo_readable = (encoder_output_fifo_level0 != 1'd0);
assign encoder_streamer_fifo_sink_valid = encoder_streamer_sink_sink_valid;
assign encoder_streamer_sink_sink_ready = encoder_streamer_fifo_sink_ready;
assign encoder_streamer_fifo_sink_first = encoder_streamer_sink_sink_first;
assign encoder_streamer_fifo_sink_last = encoder_streamer_sink_sink_last;
assign encoder_streamer_fifo_sink_payload_data = encoder_streamer_sink_sink_payload_data;
assign encoder_streamer_fifo_asyncfifo_din = {encoder_streamer_fifo_fifo_in_last, encoder_streamer_fifo_fifo_in_first, encoder_streamer_fifo_fifo_in_payload_data};
assign {encoder_streamer_fifo_fifo_out_last, encoder_streamer_fifo_fifo_out_first, encoder_streamer_fifo_fifo_out_payload_data} = encoder_streamer_fifo_asyncfifo_dout;
assign encoder_streamer_fifo_sink_ready = encoder_streamer_fifo_asyncfifo_writable;
assign encoder_streamer_fifo_asyncfifo_we = encoder_streamer_fifo_sink_valid;
assign encoder_streamer_fifo_fifo_in_first = encoder_streamer_fifo_sink_first;
assign encoder_streamer_fifo_fifo_in_last = encoder_streamer_fifo_sink_last;
assign encoder_streamer_fifo_fifo_in_payload_data = encoder_streamer_fifo_sink_payload_data;
assign encoder_streamer_fifo_source_valid = encoder_streamer_fifo_asyncfifo_readable;
assign encoder_streamer_fifo_source_first = encoder_streamer_fifo_fifo_out_first;
assign encoder_streamer_fifo_source_last = encoder_streamer_fifo_fifo_out_last;
assign encoder_streamer_fifo_source_payload_data = encoder_streamer_fifo_fifo_out_payload_data;
assign encoder_streamer_fifo_asyncfifo_re = encoder_streamer_fifo_source_ready;
assign encoder_streamer_fifo_graycounter0_ce = (encoder_streamer_fifo_asyncfifo_writable & encoder_streamer_fifo_asyncfifo_we);
assign encoder_streamer_fifo_graycounter1_ce = (encoder_streamer_fifo_asyncfifo_readable & encoder_streamer_fifo_asyncfifo_re);
assign encoder_streamer_fifo_asyncfifo_writable = (((encoder_streamer_fifo_graycounter0_q[2] == encoder_streamer_fifo_consume_wdomain[2]) | (encoder_streamer_fifo_graycounter0_q[1] == encoder_streamer_fifo_consume_wdomain[1])) | (encoder_streamer_fifo_graycounter0_q[0] != encoder_streamer_fifo_consume_wdomain[0]));
assign encoder_streamer_fifo_asyncfifo_readable = (encoder_streamer_fifo_graycounter1_q != encoder_streamer_fifo_produce_rdomain);
assign encoder_streamer_fifo_wrport_adr = encoder_streamer_fifo_graycounter0_q_binary[1:0];
assign encoder_streamer_fifo_wrport_dat_w = encoder_streamer_fifo_asyncfifo_din;
assign encoder_streamer_fifo_wrport_we = encoder_streamer_fifo_graycounter0_ce;
assign encoder_streamer_fifo_rdport_adr = encoder_streamer_fifo_graycounter1_q_next_binary[1:0];
assign encoder_streamer_fifo_asyncfifo_dout = encoder_streamer_fifo_rdport_dat_r;

// synthesis translate_off
reg dummy_d_142;
// synthesis translate_on
always @(*) begin
	encoder_streamer_fifo_graycounter0_q_next_binary <= 3'd0;
	if (encoder_streamer_fifo_graycounter0_ce) begin
		encoder_streamer_fifo_graycounter0_q_next_binary <= (encoder_streamer_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		encoder_streamer_fifo_graycounter0_q_next_binary <= encoder_streamer_fifo_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_142 <= dummy_s;
// synthesis translate_on
end
assign encoder_streamer_fifo_graycounter0_q_next = (encoder_streamer_fifo_graycounter0_q_next_binary ^ encoder_streamer_fifo_graycounter0_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_143;
// synthesis translate_on
always @(*) begin
	encoder_streamer_fifo_graycounter1_q_next_binary <= 3'd0;
	if (encoder_streamer_fifo_graycounter1_ce) begin
		encoder_streamer_fifo_graycounter1_q_next_binary <= (encoder_streamer_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		encoder_streamer_fifo_graycounter1_q_next_binary <= encoder_streamer_fifo_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_143 <= dummy_s;
// synthesis translate_on
end
assign encoder_streamer_fifo_graycounter1_q_next = (encoder_streamer_fifo_graycounter1_q_next_binary ^ encoder_streamer_fifo_graycounter1_q_next_binary[2:1]);
assign hdmi2usbsoc_interface0_wb_sdram_adr = comb_rhs_array_muxed40;
assign hdmi2usbsoc_interface0_wb_sdram_dat_w = comb_rhs_array_muxed41;
assign hdmi2usbsoc_interface0_wb_sdram_sel = comb_rhs_array_muxed42;
assign hdmi2usbsoc_interface0_wb_sdram_cyc = comb_rhs_array_muxed43;
assign hdmi2usbsoc_interface0_wb_sdram_stb = comb_rhs_array_muxed44;
assign hdmi2usbsoc_interface0_wb_sdram_we = comb_rhs_array_muxed45;
assign hdmi2usbsoc_interface0_wb_sdram_cti = comb_rhs_array_muxed46;
assign hdmi2usbsoc_interface0_wb_sdram_bte = comb_rhs_array_muxed47;
assign hdmi2usbsoc_interface1_wb_sdram_dat_r = hdmi2usbsoc_interface0_wb_sdram_dat_r;
assign hdmi2usbsoc_interface1_wb_sdram_ack = (hdmi2usbsoc_interface0_wb_sdram_ack & (wb_sdram_con_grant == 1'd0));
assign hdmi2usbsoc_interface1_wb_sdram_err = (hdmi2usbsoc_interface0_wb_sdram_err & (wb_sdram_con_grant == 1'd0));
assign wb_sdram_con_request = {hdmi2usbsoc_interface1_wb_sdram_cyc};
assign wb_sdram_con_grant = 1'd0;
assign hdmi2usbsoc_shared_adr = comb_rhs_array_muxed48;
assign hdmi2usbsoc_shared_dat_w = comb_rhs_array_muxed49;
assign hdmi2usbsoc_shared_sel = comb_rhs_array_muxed50;
assign hdmi2usbsoc_shared_cyc = comb_rhs_array_muxed51;
assign hdmi2usbsoc_shared_stb = comb_rhs_array_muxed52;
assign hdmi2usbsoc_shared_we = comb_rhs_array_muxed53;
assign hdmi2usbsoc_shared_cti = comb_rhs_array_muxed54;
assign hdmi2usbsoc_shared_bte = comb_rhs_array_muxed55;
assign hdmi2usbsoc_hdmi2usbsoc_ibus_dat_r = hdmi2usbsoc_shared_dat_r;
assign hdmi2usbsoc_hdmi2usbsoc_dbus_dat_r = hdmi2usbsoc_shared_dat_r;
assign hdmi2usbsoc_hdmi2usbsoc_ibus_ack = (hdmi2usbsoc_shared_ack & (hdmi2usbsoc_grant == 1'd0));
assign hdmi2usbsoc_hdmi2usbsoc_dbus_ack = (hdmi2usbsoc_shared_ack & (hdmi2usbsoc_grant == 1'd1));
assign hdmi2usbsoc_hdmi2usbsoc_ibus_err = (hdmi2usbsoc_shared_err & (hdmi2usbsoc_grant == 1'd0));
assign hdmi2usbsoc_hdmi2usbsoc_dbus_err = (hdmi2usbsoc_shared_err & (hdmi2usbsoc_grant == 1'd1));
assign hdmi2usbsoc_request = {hdmi2usbsoc_hdmi2usbsoc_dbus_cyc, hdmi2usbsoc_hdmi2usbsoc_ibus_cyc};

// synthesis translate_off
reg dummy_d_144;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_slave_sel <= 6'd0;
	hdmi2usbsoc_slave_sel[0] <= (hdmi2usbsoc_shared_adr[28:26] == 1'd0);
	hdmi2usbsoc_slave_sel[1] <= (hdmi2usbsoc_shared_adr[28:26] == 1'd1);
	hdmi2usbsoc_slave_sel[2] <= (hdmi2usbsoc_shared_adr[28:26] == 3'd6);
	hdmi2usbsoc_slave_sel[3] <= (hdmi2usbsoc_shared_adr[28:26] == 2'd2);
	hdmi2usbsoc_slave_sel[4] <= (hdmi2usbsoc_shared_adr[28:26] == 3'd4);
	hdmi2usbsoc_slave_sel[5] <= (hdmi2usbsoc_shared_adr[28:26] == 3'd5);
// synthesis translate_off
	dummy_d_144 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_adr = hdmi2usbsoc_shared_adr;
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_dat_w = hdmi2usbsoc_shared_dat_w;
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_sel = hdmi2usbsoc_shared_sel;
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_stb = hdmi2usbsoc_shared_stb;
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_we = hdmi2usbsoc_shared_we;
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_cti = hdmi2usbsoc_shared_cti;
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_bte = hdmi2usbsoc_shared_bte;
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_adr = hdmi2usbsoc_shared_adr;
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_dat_w = hdmi2usbsoc_shared_dat_w;
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_sel = hdmi2usbsoc_shared_sel;
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_stb = hdmi2usbsoc_shared_stb;
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_we = hdmi2usbsoc_shared_we;
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_cti = hdmi2usbsoc_shared_cti;
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_bte = hdmi2usbsoc_shared_bte;
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_adr = hdmi2usbsoc_shared_adr;
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_dat_w = hdmi2usbsoc_shared_dat_w;
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_sel = hdmi2usbsoc_shared_sel;
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_stb = hdmi2usbsoc_shared_stb;
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_we = hdmi2usbsoc_shared_we;
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_cti = hdmi2usbsoc_shared_cti;
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_bte = hdmi2usbsoc_shared_bte;
assign hdmi2usbsoc_bus_adr = hdmi2usbsoc_shared_adr;
assign hdmi2usbsoc_bus_dat_w = hdmi2usbsoc_shared_dat_w;
assign hdmi2usbsoc_bus_sel = hdmi2usbsoc_shared_sel;
assign hdmi2usbsoc_bus_stb = hdmi2usbsoc_shared_stb;
assign hdmi2usbsoc_bus_we = hdmi2usbsoc_shared_we;
assign hdmi2usbsoc_bus_cti = hdmi2usbsoc_shared_cti;
assign hdmi2usbsoc_bus_bte = hdmi2usbsoc_shared_bte;
assign hdmi2usbsoc_interface1_wb_sdram_adr = hdmi2usbsoc_shared_adr;
assign hdmi2usbsoc_interface1_wb_sdram_dat_w = hdmi2usbsoc_shared_dat_w;
assign hdmi2usbsoc_interface1_wb_sdram_sel = hdmi2usbsoc_shared_sel;
assign hdmi2usbsoc_interface1_wb_sdram_stb = hdmi2usbsoc_shared_stb;
assign hdmi2usbsoc_interface1_wb_sdram_we = hdmi2usbsoc_shared_we;
assign hdmi2usbsoc_interface1_wb_sdram_cti = hdmi2usbsoc_shared_cti;
assign hdmi2usbsoc_interface1_wb_sdram_bte = hdmi2usbsoc_shared_bte;
assign encoder_bus_adr = hdmi2usbsoc_shared_adr;
assign encoder_bus_dat_w = hdmi2usbsoc_shared_dat_w;
assign encoder_bus_sel = hdmi2usbsoc_shared_sel;
assign encoder_bus_stb = hdmi2usbsoc_shared_stb;
assign encoder_bus_we = hdmi2usbsoc_shared_we;
assign encoder_bus_cti = hdmi2usbsoc_shared_cti;
assign encoder_bus_bte = hdmi2usbsoc_shared_bte;
assign hdmi2usbsoc_hdmi2usbsoc_rom_bus_cyc = (hdmi2usbsoc_shared_cyc & hdmi2usbsoc_slave_sel[0]);
assign hdmi2usbsoc_hdmi2usbsoc_sram_bus_cyc = (hdmi2usbsoc_shared_cyc & hdmi2usbsoc_slave_sel[1]);
assign hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_cyc = (hdmi2usbsoc_shared_cyc & hdmi2usbsoc_slave_sel[2]);
assign hdmi2usbsoc_bus_cyc = (hdmi2usbsoc_shared_cyc & hdmi2usbsoc_slave_sel[3]);
assign hdmi2usbsoc_interface1_wb_sdram_cyc = (hdmi2usbsoc_shared_cyc & hdmi2usbsoc_slave_sel[4]);
assign encoder_bus_cyc = (hdmi2usbsoc_shared_cyc & hdmi2usbsoc_slave_sel[5]);
assign hdmi2usbsoc_shared_ack = (((((hdmi2usbsoc_hdmi2usbsoc_rom_bus_ack | hdmi2usbsoc_hdmi2usbsoc_sram_bus_ack) | hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_ack) | hdmi2usbsoc_bus_ack) | hdmi2usbsoc_interface1_wb_sdram_ack) | encoder_bus_ack);
assign hdmi2usbsoc_shared_err = (((((hdmi2usbsoc_hdmi2usbsoc_rom_bus_err | hdmi2usbsoc_hdmi2usbsoc_sram_bus_err) | hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_err) | hdmi2usbsoc_bus_err) | hdmi2usbsoc_interface1_wb_sdram_err) | encoder_bus_err);
assign hdmi2usbsoc_shared_dat_r = (((((({32{hdmi2usbsoc_slave_sel_r[0]}} & hdmi2usbsoc_hdmi2usbsoc_rom_bus_dat_r) | ({32{hdmi2usbsoc_slave_sel_r[1]}} & hdmi2usbsoc_hdmi2usbsoc_sram_bus_dat_r)) | ({32{hdmi2usbsoc_slave_sel_r[2]}} & hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_dat_r)) | ({32{hdmi2usbsoc_slave_sel_r[3]}} & hdmi2usbsoc_bus_dat_r)) | ({32{hdmi2usbsoc_slave_sel_r[4]}} & hdmi2usbsoc_interface1_wb_sdram_dat_r)) | ({32{hdmi2usbsoc_slave_sel_r[5]}} & encoder_bus_dat_r));
assign hdmi2usbsoc_csrbank0_sel = (hdmi2usbsoc_interface0_bank_bus_adr[13:9] == 5'd19);
assign hdmi2usbsoc_csrbank0_base3_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_base3_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 1'd0));
assign hdmi2usbsoc_csrbank0_base2_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_base2_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 1'd1));
assign hdmi2usbsoc_csrbank0_base1_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_base1_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 2'd2));
assign hdmi2usbsoc_csrbank0_base0_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_base0_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 2'd3));
assign hdmi2usbsoc_csrbank0_h_width1_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_h_width1_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 3'd4));
assign hdmi2usbsoc_csrbank0_h_width0_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_h_width0_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 3'd5));
assign hdmi2usbsoc_csrbank0_v_width1_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_v_width1_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 3'd6));
assign hdmi2usbsoc_csrbank0_v_width0_r = hdmi2usbsoc_interface0_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank0_v_width0_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 3'd7));
assign encoder_reader_start_r = hdmi2usbsoc_interface0_bank_bus_dat_w[0];
assign encoder_reader_start_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 4'd8));
assign hdmi2usbsoc_csrbank0_done_r = hdmi2usbsoc_interface0_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank0_done_re = ((hdmi2usbsoc_csrbank0_sel & hdmi2usbsoc_interface0_bank_bus_we) & (hdmi2usbsoc_interface0_bank_bus_adr[3:0] == 4'd9));
assign encoder_reader_base_storage = encoder_reader_base_storage_full[31:0];
assign hdmi2usbsoc_csrbank0_base3_w = encoder_reader_base_storage_full[31:24];
assign hdmi2usbsoc_csrbank0_base2_w = encoder_reader_base_storage_full[23:16];
assign hdmi2usbsoc_csrbank0_base1_w = encoder_reader_base_storage_full[15:8];
assign hdmi2usbsoc_csrbank0_base0_w = encoder_reader_base_storage_full[7:0];
assign encoder_reader_h_width_storage = encoder_reader_h_width_storage_full[15:0];
assign hdmi2usbsoc_csrbank0_h_width1_w = encoder_reader_h_width_storage_full[15:8];
assign hdmi2usbsoc_csrbank0_h_width0_w = encoder_reader_h_width_storage_full[7:0];
assign encoder_reader_v_width_storage = encoder_reader_v_width_storage_full[15:0];
assign hdmi2usbsoc_csrbank0_v_width1_w = encoder_reader_v_width_storage_full[15:8];
assign hdmi2usbsoc_csrbank0_v_width0_w = encoder_reader_v_width_storage_full[7:0];
assign hdmi2usbsoc_csrbank0_done_w = encoder_reader_status;
assign hdmi2usbsoc_sram0_sel = (hdmi2usbsoc_interface0_sram_bus_adr[13:9] == 5'd16);

// synthesis translate_off
reg dummy_d_145;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_interface0_sram_bus_dat_r <= 8'd0;
	if (hdmi2usbsoc_sram0_sel_r) begin
		hdmi2usbsoc_interface0_sram_bus_dat_r <= hdmi2usbsoc_sram0_dat_r;
	end
// synthesis translate_off
	dummy_d_145 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sram0_we = (hdmi2usbsoc_sram0_sel & hdmi2usbsoc_interface0_sram_bus_we);
assign hdmi2usbsoc_sram0_dat_w = hdmi2usbsoc_interface0_sram_bus_dat_w;
assign hdmi2usbsoc_sram0_adr = hdmi2usbsoc_interface0_sram_bus_adr[6:0];
assign hdmi2usbsoc_csrbank1_sel = (hdmi2usbsoc_interface1_bank_bus_adr[13:9] == 4'd15);
assign hdmi2usbsoc_csrbank1_edid_hpd_notif_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_edid_hpd_notif_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 1'd0));
assign hdmi2usbsoc_csrbank1_edid_hpd_en0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_edid_hpd_en0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 1'd1));
assign hdmi2usbsoc_csrbank1_clocking_pll_reset0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_clocking_pll_reset0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 2'd2));
assign hdmi2usbsoc_csrbank1_clocking_locked_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_clocking_locked_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 2'd3));
assign hdmi2usbsoc_csrbank1_clocking_pll_adr0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[4:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_adr0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 3'd4));
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_r1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_r1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 3'd5));
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_r0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_r0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 3'd6));
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 3'd7));
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd8));
assign hdmi2usbsoc_hdmi_in0_pll_read_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_pll_read_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd9));
assign hdmi2usbsoc_hdmi_in0_pll_write_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_pll_write_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd10));
assign hdmi2usbsoc_csrbank1_clocking_pll_drdy_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_clocking_pll_drdy_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd11));
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_r = hdmi2usbsoc_interface1_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd12));
assign hdmi2usbsoc_csrbank1_data0_cap_dly_busy_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_data0_cap_dly_busy_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd13));
assign hdmi2usbsoc_csrbank1_data0_cap_phase_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_data0_cap_phase_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd14));
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_reset_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_reset_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 4'd15));
assign hdmi2usbsoc_csrbank1_data0_charsync_char_synced_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_data0_charsync_char_synced_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd16));
assign hdmi2usbsoc_csrbank1_data0_charsync_ctl_pos_r = hdmi2usbsoc_interface1_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank1_data0_charsync_ctl_pos_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd17));
assign hdmi2usbsoc_hdmi_in0_wer0_update_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_wer0_update_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd18));
assign hdmi2usbsoc_csrbank1_data0_wer_value2_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data0_wer_value2_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd19));
assign hdmi2usbsoc_csrbank1_data0_wer_value1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data0_wer_value1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd20));
assign hdmi2usbsoc_csrbank1_data0_wer_value0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data0_wer_value0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd21));
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_r = hdmi2usbsoc_interface1_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd22));
assign hdmi2usbsoc_csrbank1_data1_cap_dly_busy_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_data1_cap_dly_busy_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd23));
assign hdmi2usbsoc_csrbank1_data1_cap_phase_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_data1_cap_phase_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd24));
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_reset_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_reset_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd25));
assign hdmi2usbsoc_csrbank1_data1_charsync_char_synced_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_data1_charsync_char_synced_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd26));
assign hdmi2usbsoc_csrbank1_data1_charsync_ctl_pos_r = hdmi2usbsoc_interface1_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank1_data1_charsync_ctl_pos_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd27));
assign hdmi2usbsoc_hdmi_in0_wer1_update_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_wer1_update_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd28));
assign hdmi2usbsoc_csrbank1_data1_wer_value2_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data1_wer_value2_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd29));
assign hdmi2usbsoc_csrbank1_data1_wer_value1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data1_wer_value1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd30));
assign hdmi2usbsoc_csrbank1_data1_wer_value0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data1_wer_value0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 5'd31));
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_r = hdmi2usbsoc_interface1_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd32));
assign hdmi2usbsoc_csrbank1_data2_cap_dly_busy_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_data2_cap_dly_busy_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd33));
assign hdmi2usbsoc_csrbank1_data2_cap_phase_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_data2_cap_phase_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd34));
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_reset_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_reset_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd35));
assign hdmi2usbsoc_csrbank1_data2_charsync_char_synced_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_data2_charsync_char_synced_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd36));
assign hdmi2usbsoc_csrbank1_data2_charsync_ctl_pos_r = hdmi2usbsoc_interface1_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank1_data2_charsync_ctl_pos_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd37));
assign hdmi2usbsoc_hdmi_in0_wer2_update_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_wer2_update_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd38));
assign hdmi2usbsoc_csrbank1_data2_wer_value2_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data2_wer_value2_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd39));
assign hdmi2usbsoc_csrbank1_data2_wer_value1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data2_wer_value1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd40));
assign hdmi2usbsoc_csrbank1_data2_wer_value0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_data2_wer_value0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd41));
assign hdmi2usbsoc_csrbank1_chansync_channels_synced_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank1_chansync_channels_synced_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd42));
assign hdmi2usbsoc_csrbank1_resdetection_hres1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank1_resdetection_hres1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd43));
assign hdmi2usbsoc_csrbank1_resdetection_hres0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_resdetection_hres0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd44));
assign hdmi2usbsoc_csrbank1_resdetection_vres1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank1_resdetection_vres1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd45));
assign hdmi2usbsoc_csrbank1_resdetection_vres0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_resdetection_vres0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd46));
assign hdmi2usbsoc_hdmi_in0_frame_overflow_r = hdmi2usbsoc_interface1_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in0_frame_overflow_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd47));
assign hdmi2usbsoc_csrbank1_dma_frame_size3_r = hdmi2usbsoc_interface1_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank1_dma_frame_size3_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd48));
assign hdmi2usbsoc_csrbank1_dma_frame_size2_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_frame_size2_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd49));
assign hdmi2usbsoc_csrbank1_dma_frame_size1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_frame_size1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd50));
assign hdmi2usbsoc_csrbank1_dma_frame_size0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_frame_size0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd51));
assign hdmi2usbsoc_csrbank1_dma_slot0_status0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_dma_slot0_status0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd52));
assign hdmi2usbsoc_csrbank1_dma_slot0_address3_r = hdmi2usbsoc_interface1_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank1_dma_slot0_address3_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd53));
assign hdmi2usbsoc_csrbank1_dma_slot0_address2_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_slot0_address2_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd54));
assign hdmi2usbsoc_csrbank1_dma_slot0_address1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_slot0_address1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd55));
assign hdmi2usbsoc_csrbank1_dma_slot0_address0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_slot0_address0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd56));
assign hdmi2usbsoc_csrbank1_dma_slot1_status0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_dma_slot1_status0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd57));
assign hdmi2usbsoc_csrbank1_dma_slot1_address3_r = hdmi2usbsoc_interface1_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank1_dma_slot1_address3_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd58));
assign hdmi2usbsoc_csrbank1_dma_slot1_address2_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_slot1_address2_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd59));
assign hdmi2usbsoc_csrbank1_dma_slot1_address1_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_slot1_address1_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd60));
assign hdmi2usbsoc_csrbank1_dma_slot1_address0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank1_dma_slot1_address0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd61));
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_status_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_status_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd62));
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 6'd63));
assign hdmi2usbsoc_csrbank1_dma_ev_enable0_r = hdmi2usbsoc_interface1_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank1_dma_ev_enable0_re = ((hdmi2usbsoc_csrbank1_sel & hdmi2usbsoc_interface1_bank_bus_we) & (hdmi2usbsoc_interface1_bank_bus_adr[6:0] == 7'd64));
assign hdmi2usbsoc_csrbank1_edid_hpd_notif_w = hdmi2usbsoc_hdmi_in0_edid_status;
assign hdmi2usbsoc_hdmi_in0_edid_storage = hdmi2usbsoc_hdmi_in0_edid_storage_full;
assign hdmi2usbsoc_csrbank1_edid_hpd_en0_w = hdmi2usbsoc_hdmi_in0_edid_storage_full;
assign hdmi2usbsoc_hdmi_in0_pll_reset_storage = hdmi2usbsoc_hdmi_in0_pll_reset_storage_full;
assign hdmi2usbsoc_csrbank1_clocking_pll_reset0_w = hdmi2usbsoc_hdmi_in0_pll_reset_storage_full;
assign hdmi2usbsoc_csrbank1_clocking_locked_w = hdmi2usbsoc_hdmi_in0_locked_status;
assign hdmi2usbsoc_hdmi_in0_pll_adr_storage = hdmi2usbsoc_hdmi_in0_pll_adr_storage_full[4:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_adr0_w = hdmi2usbsoc_hdmi_in0_pll_adr_storage_full[4:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_r1_w = hdmi2usbsoc_hdmi_in0_pll_dat_r_status[15:8];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_r0_w = hdmi2usbsoc_hdmi_in0_pll_dat_r_status[7:0];
assign hdmi2usbsoc_hdmi_in0_pll_dat_w_storage = hdmi2usbsoc_hdmi_in0_pll_dat_w_storage_full[15:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_w = hdmi2usbsoc_hdmi_in0_pll_dat_w_storage_full[15:8];
assign hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_w = hdmi2usbsoc_hdmi_in0_pll_dat_w_storage_full[7:0];
assign hdmi2usbsoc_csrbank1_clocking_pll_drdy_w = hdmi2usbsoc_hdmi_in0_pll_drdy_status;
assign hdmi2usbsoc_csrbank1_data0_cap_dly_busy_w = hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_busy_status[1:0];
assign hdmi2usbsoc_csrbank1_data0_cap_phase_w = hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_status[1:0];
assign hdmi2usbsoc_csrbank1_data0_charsync_char_synced_w = hdmi2usbsoc_hdmi_in0_charsync0_char_synced_status;
assign hdmi2usbsoc_csrbank1_data0_charsync_ctl_pos_w = hdmi2usbsoc_hdmi_in0_charsync0_ctl_pos_status[3:0];
assign hdmi2usbsoc_csrbank1_data0_wer_value2_w = hdmi2usbsoc_hdmi_in0_wer0_status[23:16];
assign hdmi2usbsoc_csrbank1_data0_wer_value1_w = hdmi2usbsoc_hdmi_in0_wer0_status[15:8];
assign hdmi2usbsoc_csrbank1_data0_wer_value0_w = hdmi2usbsoc_hdmi_in0_wer0_status[7:0];
assign hdmi2usbsoc_csrbank1_data1_cap_dly_busy_w = hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_busy_status[1:0];
assign hdmi2usbsoc_csrbank1_data1_cap_phase_w = hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_status[1:0];
assign hdmi2usbsoc_csrbank1_data1_charsync_char_synced_w = hdmi2usbsoc_hdmi_in0_charsync1_char_synced_status;
assign hdmi2usbsoc_csrbank1_data1_charsync_ctl_pos_w = hdmi2usbsoc_hdmi_in0_charsync1_ctl_pos_status[3:0];
assign hdmi2usbsoc_csrbank1_data1_wer_value2_w = hdmi2usbsoc_hdmi_in0_wer1_status[23:16];
assign hdmi2usbsoc_csrbank1_data1_wer_value1_w = hdmi2usbsoc_hdmi_in0_wer1_status[15:8];
assign hdmi2usbsoc_csrbank1_data1_wer_value0_w = hdmi2usbsoc_hdmi_in0_wer1_status[7:0];
assign hdmi2usbsoc_csrbank1_data2_cap_dly_busy_w = hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_busy_status[1:0];
assign hdmi2usbsoc_csrbank1_data2_cap_phase_w = hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_status[1:0];
assign hdmi2usbsoc_csrbank1_data2_charsync_char_synced_w = hdmi2usbsoc_hdmi_in0_charsync2_char_synced_status;
assign hdmi2usbsoc_csrbank1_data2_charsync_ctl_pos_w = hdmi2usbsoc_hdmi_in0_charsync2_ctl_pos_status[3:0];
assign hdmi2usbsoc_csrbank1_data2_wer_value2_w = hdmi2usbsoc_hdmi_in0_wer2_status[23:16];
assign hdmi2usbsoc_csrbank1_data2_wer_value1_w = hdmi2usbsoc_hdmi_in0_wer2_status[15:8];
assign hdmi2usbsoc_csrbank1_data2_wer_value0_w = hdmi2usbsoc_hdmi_in0_wer2_status[7:0];
assign hdmi2usbsoc_csrbank1_chansync_channels_synced_w = hdmi2usbsoc_hdmi_in0_chansync_status;
assign hdmi2usbsoc_csrbank1_resdetection_hres1_w = hdmi2usbsoc_hdmi_in0_resdetection_hres_status[10:8];
assign hdmi2usbsoc_csrbank1_resdetection_hres0_w = hdmi2usbsoc_hdmi_in0_resdetection_hres_status[7:0];
assign hdmi2usbsoc_csrbank1_resdetection_vres1_w = hdmi2usbsoc_hdmi_in0_resdetection_vres_status[10:8];
assign hdmi2usbsoc_csrbank1_resdetection_vres0_w = hdmi2usbsoc_hdmi_in0_resdetection_vres_status[7:0];
assign hdmi2usbsoc_hdmi_in0_dma_frame_size_storage = hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[26:3];
assign hdmi2usbsoc_csrbank1_dma_frame_size3_w = hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[26:24];
assign hdmi2usbsoc_csrbank1_dma_frame_size2_w = hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[23:16];
assign hdmi2usbsoc_csrbank1_dma_frame_size1_w = hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[15:8];
assign hdmi2usbsoc_csrbank1_dma_frame_size0_w = {hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[7:3], {5{1'd0}}};
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage_full[1:0];
assign hdmi2usbsoc_csrbank1_dma_slot0_status0_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage_full[1:0];
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[26:3];
assign hdmi2usbsoc_csrbank1_dma_slot0_address3_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[26:24];
assign hdmi2usbsoc_csrbank1_dma_slot0_address2_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[23:16];
assign hdmi2usbsoc_csrbank1_dma_slot0_address1_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[15:8];
assign hdmi2usbsoc_csrbank1_dma_slot0_address0_w = {hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[7:3], {5{1'd0}}};
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage_full[1:0];
assign hdmi2usbsoc_csrbank1_dma_slot1_status0_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage_full[1:0];
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[26:3];
assign hdmi2usbsoc_csrbank1_dma_slot1_address3_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[26:24];
assign hdmi2usbsoc_csrbank1_dma_slot1_address2_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[23:16];
assign hdmi2usbsoc_csrbank1_dma_slot1_address1_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[15:8];
assign hdmi2usbsoc_csrbank1_dma_slot1_address0_w = {hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[7:3], {5{1'd0}}};
assign hdmi2usbsoc_hdmi_in0_dma_slot_array_storage = hdmi2usbsoc_hdmi_in0_dma_slot_array_storage_full[1:0];
assign hdmi2usbsoc_csrbank1_dma_ev_enable0_w = hdmi2usbsoc_hdmi_in0_dma_slot_array_storage_full[1:0];
assign hdmi2usbsoc_sram1_sel = (hdmi2usbsoc_interface1_sram_bus_adr[13:9] == 5'd18);

// synthesis translate_off
reg dummy_d_146;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_interface1_sram_bus_dat_r <= 8'd0;
	if (hdmi2usbsoc_sram1_sel_r) begin
		hdmi2usbsoc_interface1_sram_bus_dat_r <= hdmi2usbsoc_sram1_dat_r;
	end
// synthesis translate_off
	dummy_d_146 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sram1_we = (hdmi2usbsoc_sram1_sel & hdmi2usbsoc_interface1_sram_bus_we);
assign hdmi2usbsoc_sram1_dat_w = hdmi2usbsoc_interface1_sram_bus_dat_w;
assign hdmi2usbsoc_sram1_adr = hdmi2usbsoc_interface1_sram_bus_adr[6:0];
assign hdmi2usbsoc_csrbank2_sel = (hdmi2usbsoc_interface2_bank_bus_adr[13:9] == 5'd17);
assign hdmi2usbsoc_csrbank2_edid_hpd_notif_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_edid_hpd_notif_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 1'd0));
assign hdmi2usbsoc_csrbank2_edid_hpd_en0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_edid_hpd_en0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 1'd1));
assign hdmi2usbsoc_csrbank2_clocking_pll_reset0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_clocking_pll_reset0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 2'd2));
assign hdmi2usbsoc_csrbank2_clocking_locked_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_clocking_locked_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 2'd3));
assign hdmi2usbsoc_csrbank2_clocking_pll_adr0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[4:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_adr0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 3'd4));
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_r1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_r1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 3'd5));
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_r0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_r0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 3'd6));
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 3'd7));
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd8));
assign hdmi2usbsoc_hdmi_in1_pll_read_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_pll_read_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd9));
assign hdmi2usbsoc_hdmi_in1_pll_write_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_pll_write_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd10));
assign hdmi2usbsoc_csrbank2_clocking_pll_drdy_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_clocking_pll_drdy_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd11));
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_r = hdmi2usbsoc_interface2_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd12));
assign hdmi2usbsoc_csrbank2_data0_cap_dly_busy_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_data0_cap_dly_busy_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd13));
assign hdmi2usbsoc_csrbank2_data0_cap_phase_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_data0_cap_phase_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd14));
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_reset_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_reset_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 4'd15));
assign hdmi2usbsoc_csrbank2_data0_charsync_char_synced_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_data0_charsync_char_synced_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd16));
assign hdmi2usbsoc_csrbank2_data0_charsync_ctl_pos_r = hdmi2usbsoc_interface2_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank2_data0_charsync_ctl_pos_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd17));
assign hdmi2usbsoc_hdmi_in1_wer0_update_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_wer0_update_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd18));
assign hdmi2usbsoc_csrbank2_data0_wer_value2_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data0_wer_value2_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd19));
assign hdmi2usbsoc_csrbank2_data0_wer_value1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data0_wer_value1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd20));
assign hdmi2usbsoc_csrbank2_data0_wer_value0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data0_wer_value0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd21));
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_r = hdmi2usbsoc_interface2_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd22));
assign hdmi2usbsoc_csrbank2_data1_cap_dly_busy_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_data1_cap_dly_busy_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd23));
assign hdmi2usbsoc_csrbank2_data1_cap_phase_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_data1_cap_phase_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd24));
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_reset_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_reset_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd25));
assign hdmi2usbsoc_csrbank2_data1_charsync_char_synced_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_data1_charsync_char_synced_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd26));
assign hdmi2usbsoc_csrbank2_data1_charsync_ctl_pos_r = hdmi2usbsoc_interface2_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank2_data1_charsync_ctl_pos_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd27));
assign hdmi2usbsoc_hdmi_in1_wer1_update_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_wer1_update_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd28));
assign hdmi2usbsoc_csrbank2_data1_wer_value2_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data1_wer_value2_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd29));
assign hdmi2usbsoc_csrbank2_data1_wer_value1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data1_wer_value1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd30));
assign hdmi2usbsoc_csrbank2_data1_wer_value0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data1_wer_value0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 5'd31));
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_r = hdmi2usbsoc_interface2_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd32));
assign hdmi2usbsoc_csrbank2_data2_cap_dly_busy_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_data2_cap_dly_busy_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd33));
assign hdmi2usbsoc_csrbank2_data2_cap_phase_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_data2_cap_phase_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd34));
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_reset_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_reset_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd35));
assign hdmi2usbsoc_csrbank2_data2_charsync_char_synced_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_data2_charsync_char_synced_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd36));
assign hdmi2usbsoc_csrbank2_data2_charsync_ctl_pos_r = hdmi2usbsoc_interface2_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank2_data2_charsync_ctl_pos_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd37));
assign hdmi2usbsoc_hdmi_in1_wer2_update_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_wer2_update_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd38));
assign hdmi2usbsoc_csrbank2_data2_wer_value2_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data2_wer_value2_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd39));
assign hdmi2usbsoc_csrbank2_data2_wer_value1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data2_wer_value1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd40));
assign hdmi2usbsoc_csrbank2_data2_wer_value0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_data2_wer_value0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd41));
assign hdmi2usbsoc_csrbank2_chansync_channels_synced_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank2_chansync_channels_synced_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd42));
assign hdmi2usbsoc_csrbank2_resdetection_hres1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank2_resdetection_hres1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd43));
assign hdmi2usbsoc_csrbank2_resdetection_hres0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_resdetection_hres0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd44));
assign hdmi2usbsoc_csrbank2_resdetection_vres1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank2_resdetection_vres1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd45));
assign hdmi2usbsoc_csrbank2_resdetection_vres0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_resdetection_vres0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd46));
assign hdmi2usbsoc_hdmi_in1_frame_overflow_r = hdmi2usbsoc_interface2_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_in1_frame_overflow_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd47));
assign hdmi2usbsoc_csrbank2_dma_frame_size3_r = hdmi2usbsoc_interface2_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank2_dma_frame_size3_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd48));
assign hdmi2usbsoc_csrbank2_dma_frame_size2_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_frame_size2_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd49));
assign hdmi2usbsoc_csrbank2_dma_frame_size1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_frame_size1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd50));
assign hdmi2usbsoc_csrbank2_dma_frame_size0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_frame_size0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd51));
assign hdmi2usbsoc_csrbank2_dma_slot0_status0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_dma_slot0_status0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd52));
assign hdmi2usbsoc_csrbank2_dma_slot0_address3_r = hdmi2usbsoc_interface2_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank2_dma_slot0_address3_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd53));
assign hdmi2usbsoc_csrbank2_dma_slot0_address2_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_slot0_address2_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd54));
assign hdmi2usbsoc_csrbank2_dma_slot0_address1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_slot0_address1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd55));
assign hdmi2usbsoc_csrbank2_dma_slot0_address0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_slot0_address0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd56));
assign hdmi2usbsoc_csrbank2_dma_slot1_status0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_dma_slot1_status0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd57));
assign hdmi2usbsoc_csrbank2_dma_slot1_address3_r = hdmi2usbsoc_interface2_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank2_dma_slot1_address3_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd58));
assign hdmi2usbsoc_csrbank2_dma_slot1_address2_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_slot1_address2_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd59));
assign hdmi2usbsoc_csrbank2_dma_slot1_address1_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_slot1_address1_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd60));
assign hdmi2usbsoc_csrbank2_dma_slot1_address0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank2_dma_slot1_address0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd61));
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_status_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_status_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd62));
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 6'd63));
assign hdmi2usbsoc_csrbank2_dma_ev_enable0_r = hdmi2usbsoc_interface2_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank2_dma_ev_enable0_re = ((hdmi2usbsoc_csrbank2_sel & hdmi2usbsoc_interface2_bank_bus_we) & (hdmi2usbsoc_interface2_bank_bus_adr[6:0] == 7'd64));
assign hdmi2usbsoc_csrbank2_edid_hpd_notif_w = hdmi2usbsoc_hdmi_in1_edid_status;
assign hdmi2usbsoc_hdmi_in1_edid_storage = hdmi2usbsoc_hdmi_in1_edid_storage_full;
assign hdmi2usbsoc_csrbank2_edid_hpd_en0_w = hdmi2usbsoc_hdmi_in1_edid_storage_full;
assign hdmi2usbsoc_hdmi_in1_pll_reset_storage = hdmi2usbsoc_hdmi_in1_pll_reset_storage_full;
assign hdmi2usbsoc_csrbank2_clocking_pll_reset0_w = hdmi2usbsoc_hdmi_in1_pll_reset_storage_full;
assign hdmi2usbsoc_csrbank2_clocking_locked_w = hdmi2usbsoc_hdmi_in1_locked_status;
assign hdmi2usbsoc_hdmi_in1_pll_adr_storage = hdmi2usbsoc_hdmi_in1_pll_adr_storage_full[4:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_adr0_w = hdmi2usbsoc_hdmi_in1_pll_adr_storage_full[4:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_r1_w = hdmi2usbsoc_hdmi_in1_pll_dat_r_status[15:8];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_r0_w = hdmi2usbsoc_hdmi_in1_pll_dat_r_status[7:0];
assign hdmi2usbsoc_hdmi_in1_pll_dat_w_storage = hdmi2usbsoc_hdmi_in1_pll_dat_w_storage_full[15:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_w = hdmi2usbsoc_hdmi_in1_pll_dat_w_storage_full[15:8];
assign hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_w = hdmi2usbsoc_hdmi_in1_pll_dat_w_storage_full[7:0];
assign hdmi2usbsoc_csrbank2_clocking_pll_drdy_w = hdmi2usbsoc_hdmi_in1_pll_drdy_status;
assign hdmi2usbsoc_csrbank2_data0_cap_dly_busy_w = hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_busy_status[1:0];
assign hdmi2usbsoc_csrbank2_data0_cap_phase_w = hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_status[1:0];
assign hdmi2usbsoc_csrbank2_data0_charsync_char_synced_w = hdmi2usbsoc_hdmi_in1_charsync0_char_synced_status;
assign hdmi2usbsoc_csrbank2_data0_charsync_ctl_pos_w = hdmi2usbsoc_hdmi_in1_charsync0_ctl_pos_status[3:0];
assign hdmi2usbsoc_csrbank2_data0_wer_value2_w = hdmi2usbsoc_hdmi_in1_wer0_status[23:16];
assign hdmi2usbsoc_csrbank2_data0_wer_value1_w = hdmi2usbsoc_hdmi_in1_wer0_status[15:8];
assign hdmi2usbsoc_csrbank2_data0_wer_value0_w = hdmi2usbsoc_hdmi_in1_wer0_status[7:0];
assign hdmi2usbsoc_csrbank2_data1_cap_dly_busy_w = hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_busy_status[1:0];
assign hdmi2usbsoc_csrbank2_data1_cap_phase_w = hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_status[1:0];
assign hdmi2usbsoc_csrbank2_data1_charsync_char_synced_w = hdmi2usbsoc_hdmi_in1_charsync1_char_synced_status;
assign hdmi2usbsoc_csrbank2_data1_charsync_ctl_pos_w = hdmi2usbsoc_hdmi_in1_charsync1_ctl_pos_status[3:0];
assign hdmi2usbsoc_csrbank2_data1_wer_value2_w = hdmi2usbsoc_hdmi_in1_wer1_status[23:16];
assign hdmi2usbsoc_csrbank2_data1_wer_value1_w = hdmi2usbsoc_hdmi_in1_wer1_status[15:8];
assign hdmi2usbsoc_csrbank2_data1_wer_value0_w = hdmi2usbsoc_hdmi_in1_wer1_status[7:0];
assign hdmi2usbsoc_csrbank2_data2_cap_dly_busy_w = hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_busy_status[1:0];
assign hdmi2usbsoc_csrbank2_data2_cap_phase_w = hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_status[1:0];
assign hdmi2usbsoc_csrbank2_data2_charsync_char_synced_w = hdmi2usbsoc_hdmi_in1_charsync2_char_synced_status;
assign hdmi2usbsoc_csrbank2_data2_charsync_ctl_pos_w = hdmi2usbsoc_hdmi_in1_charsync2_ctl_pos_status[3:0];
assign hdmi2usbsoc_csrbank2_data2_wer_value2_w = hdmi2usbsoc_hdmi_in1_wer2_status[23:16];
assign hdmi2usbsoc_csrbank2_data2_wer_value1_w = hdmi2usbsoc_hdmi_in1_wer2_status[15:8];
assign hdmi2usbsoc_csrbank2_data2_wer_value0_w = hdmi2usbsoc_hdmi_in1_wer2_status[7:0];
assign hdmi2usbsoc_csrbank2_chansync_channels_synced_w = hdmi2usbsoc_hdmi_in1_chansync_status;
assign hdmi2usbsoc_csrbank2_resdetection_hres1_w = hdmi2usbsoc_hdmi_in1_resdetection_hres_status[10:8];
assign hdmi2usbsoc_csrbank2_resdetection_hres0_w = hdmi2usbsoc_hdmi_in1_resdetection_hres_status[7:0];
assign hdmi2usbsoc_csrbank2_resdetection_vres1_w = hdmi2usbsoc_hdmi_in1_resdetection_vres_status[10:8];
assign hdmi2usbsoc_csrbank2_resdetection_vres0_w = hdmi2usbsoc_hdmi_in1_resdetection_vres_status[7:0];
assign hdmi2usbsoc_hdmi_in1_dma_frame_size_storage = hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[26:3];
assign hdmi2usbsoc_csrbank2_dma_frame_size3_w = hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[26:24];
assign hdmi2usbsoc_csrbank2_dma_frame_size2_w = hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[23:16];
assign hdmi2usbsoc_csrbank2_dma_frame_size1_w = hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[15:8];
assign hdmi2usbsoc_csrbank2_dma_frame_size0_w = {hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[7:3], {5{1'd0}}};
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage_full[1:0];
assign hdmi2usbsoc_csrbank2_dma_slot0_status0_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage_full[1:0];
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[26:3];
assign hdmi2usbsoc_csrbank2_dma_slot0_address3_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[26:24];
assign hdmi2usbsoc_csrbank2_dma_slot0_address2_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[23:16];
assign hdmi2usbsoc_csrbank2_dma_slot0_address1_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[15:8];
assign hdmi2usbsoc_csrbank2_dma_slot0_address0_w = {hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[7:3], {5{1'd0}}};
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage_full[1:0];
assign hdmi2usbsoc_csrbank2_dma_slot1_status0_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage_full[1:0];
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[26:3];
assign hdmi2usbsoc_csrbank2_dma_slot1_address3_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[26:24];
assign hdmi2usbsoc_csrbank2_dma_slot1_address2_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[23:16];
assign hdmi2usbsoc_csrbank2_dma_slot1_address1_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[15:8];
assign hdmi2usbsoc_csrbank2_dma_slot1_address0_w = {hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[7:3], {5{1'd0}}};
assign hdmi2usbsoc_hdmi_in1_dma_slot_array_storage = hdmi2usbsoc_hdmi_in1_dma_slot_array_storage_full[1:0];
assign hdmi2usbsoc_csrbank2_dma_ev_enable0_w = hdmi2usbsoc_hdmi_in1_dma_slot_array_storage_full[1:0];
assign hdmi2usbsoc_csrbank3_sel = (hdmi2usbsoc_interface3_bank_bus_adr[13:9] == 4'd13);
assign hdmi2usbsoc_csrbank3_core_underflow_enable0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank3_core_underflow_enable0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 1'd0));
assign hdmi2usbsoc_hdmi_out0_core_underflow_update_underflow_update_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_out0_core_underflow_update_underflow_update_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 1'd1));
assign hdmi2usbsoc_csrbank3_core_underflow_counter3_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_underflow_counter3_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 2'd2));
assign hdmi2usbsoc_csrbank3_core_underflow_counter2_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_underflow_counter2_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 2'd3));
assign hdmi2usbsoc_csrbank3_core_underflow_counter1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_underflow_counter1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 3'd4));
assign hdmi2usbsoc_csrbank3_core_underflow_counter0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_underflow_counter0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 3'd5));
assign hdmi2usbsoc_csrbank3_core_initiator_enable0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank3_core_initiator_enable0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 3'd6));
assign hdmi2usbsoc_csrbank3_core_initiator_hres1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hres1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 3'd7));
assign hdmi2usbsoc_csrbank3_core_initiator_hres0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hres0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd8));
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd9));
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd10));
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd11));
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd12));
assign hdmi2usbsoc_csrbank3_core_initiator_hscan1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hscan1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd13));
assign hdmi2usbsoc_csrbank3_core_initiator_hscan0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hscan0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd14));
assign hdmi2usbsoc_csrbank3_core_initiator_vres1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vres1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 4'd15));
assign hdmi2usbsoc_csrbank3_core_initiator_vres0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vres0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd16));
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd17));
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd18));
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd19));
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd20));
assign hdmi2usbsoc_csrbank3_core_initiator_vscan1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vscan1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd21));
assign hdmi2usbsoc_csrbank3_core_initiator_vscan0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vscan0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd22));
assign hdmi2usbsoc_csrbank3_core_initiator_base3_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_base3_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd23));
assign hdmi2usbsoc_csrbank3_core_initiator_base2_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_base2_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd24));
assign hdmi2usbsoc_csrbank3_core_initiator_base1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_base1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd25));
assign hdmi2usbsoc_csrbank3_core_initiator_base0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_base0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd26));
assign hdmi2usbsoc_csrbank3_core_initiator_length3_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_length3_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd27));
assign hdmi2usbsoc_csrbank3_core_initiator_length2_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_length2_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd28));
assign hdmi2usbsoc_csrbank3_core_initiator_length1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_length1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd29));
assign hdmi2usbsoc_csrbank3_core_initiator_length0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_core_initiator_length0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd30));
assign hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 5'd31));
assign hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd32));
assign hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd33));
assign hdmi2usbsoc_hdmi_out0_driver_clocking_send_go_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_out0_driver_clocking_send_go_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd34));
assign hdmi2usbsoc_csrbank3_driver_clocking_status_r = hdmi2usbsoc_interface3_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_status_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd35));
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd36));
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[4:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd37));
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd38));
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd39));
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd40));
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_r = hdmi2usbsoc_interface3_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd41));
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd42));
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd43));
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_drdy_r = hdmi2usbsoc_interface3_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_drdy_re = ((hdmi2usbsoc_csrbank3_sel & hdmi2usbsoc_interface3_bank_bus_we) & (hdmi2usbsoc_interface3_bank_bus_adr[5:0] == 6'd44));
assign hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage = hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage_full;
assign hdmi2usbsoc_csrbank3_core_underflow_enable0_w = hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage_full;
assign hdmi2usbsoc_csrbank3_core_underflow_counter3_w = hdmi2usbsoc_hdmi_out0_core_underflow_counter_status[31:24];
assign hdmi2usbsoc_csrbank3_core_underflow_counter2_w = hdmi2usbsoc_hdmi_out0_core_underflow_counter_status[23:16];
assign hdmi2usbsoc_csrbank3_core_underflow_counter1_w = hdmi2usbsoc_hdmi_out0_core_underflow_counter_status[15:8];
assign hdmi2usbsoc_csrbank3_core_underflow_counter0_w = hdmi2usbsoc_hdmi_out0_core_underflow_counter_status[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage = hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage_full;
assign hdmi2usbsoc_csrbank3_core_initiator_enable0_w = hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage_full;
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hres1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_hres0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_hscan1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_hscan0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vres1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_vres0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage_full[11:0];
assign hdmi2usbsoc_csrbank3_core_initiator_vscan1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage_full[11:8];
assign hdmi2usbsoc_csrbank3_core_initiator_vscan0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full[31:0];
assign hdmi2usbsoc_csrbank3_core_initiator_base3_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full[31:24];
assign hdmi2usbsoc_csrbank3_core_initiator_base2_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full[23:16];
assign hdmi2usbsoc_csrbank3_core_initiator_base1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full[15:8];
assign hdmi2usbsoc_csrbank3_core_initiator_base0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full[31:0];
assign hdmi2usbsoc_csrbank3_core_initiator_length3_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full[31:24];
assign hdmi2usbsoc_csrbank3_core_initiator_length2_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full[23:16];
assign hdmi2usbsoc_csrbank3_core_initiator_length1_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full[15:8];
assign hdmi2usbsoc_csrbank3_core_initiator_length0_w = hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage = hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage_full[9:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_w = hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage_full[9:8];
assign hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_w = hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage_full[7:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_status_w = hdmi2usbsoc_hdmi_out0_driver_clocking_status_status[3:0];
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage_full;
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_w = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage_full;
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage_full[4:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_w = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage_full[4:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r1_w = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_r_status[15:8];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r0_w = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_r_status[7:0];
assign hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage_full[15:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_w = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage_full[15:8];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_w = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage_full[7:0];
assign hdmi2usbsoc_csrbank3_driver_clocking_pll_drdy_w = hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy_status;
assign hdmi2usbsoc_csrbank4_sel = (hdmi2usbsoc_interface4_bank_bus_adr[13:9] == 4'd14);
assign hdmi2usbsoc_csrbank4_core_underflow_enable0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank4_core_underflow_enable0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 1'd0));
assign hdmi2usbsoc_hdmi_out1_core_underflow_update_underflow_update_r = hdmi2usbsoc_interface4_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi_out1_core_underflow_update_underflow_update_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 1'd1));
assign hdmi2usbsoc_csrbank4_core_underflow_counter3_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_underflow_counter3_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 2'd2));
assign hdmi2usbsoc_csrbank4_core_underflow_counter2_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_underflow_counter2_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 2'd3));
assign hdmi2usbsoc_csrbank4_core_underflow_counter1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_underflow_counter1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 3'd4));
assign hdmi2usbsoc_csrbank4_core_underflow_counter0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_underflow_counter0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 3'd5));
assign hdmi2usbsoc_csrbank4_core_initiator_enable0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank4_core_initiator_enable0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 3'd6));
assign hdmi2usbsoc_csrbank4_core_initiator_hres1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hres1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 3'd7));
assign hdmi2usbsoc_csrbank4_core_initiator_hres0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hres0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd8));
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd9));
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd10));
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd11));
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd12));
assign hdmi2usbsoc_csrbank4_core_initiator_hscan1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hscan1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd13));
assign hdmi2usbsoc_csrbank4_core_initiator_hscan0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hscan0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd14));
assign hdmi2usbsoc_csrbank4_core_initiator_vres1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vres1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 4'd15));
assign hdmi2usbsoc_csrbank4_core_initiator_vres0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vres0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd16));
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd17));
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd18));
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd19));
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd20));
assign hdmi2usbsoc_csrbank4_core_initiator_vscan1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vscan1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd21));
assign hdmi2usbsoc_csrbank4_core_initiator_vscan0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vscan0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd22));
assign hdmi2usbsoc_csrbank4_core_initiator_base3_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_base3_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd23));
assign hdmi2usbsoc_csrbank4_core_initiator_base2_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_base2_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd24));
assign hdmi2usbsoc_csrbank4_core_initiator_base1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_base1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd25));
assign hdmi2usbsoc_csrbank4_core_initiator_base0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_base0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd26));
assign hdmi2usbsoc_csrbank4_core_initiator_length3_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_length3_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd27));
assign hdmi2usbsoc_csrbank4_core_initiator_length2_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_length2_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd28));
assign hdmi2usbsoc_csrbank4_core_initiator_length1_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_length1_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd29));
assign hdmi2usbsoc_csrbank4_core_initiator_length0_r = hdmi2usbsoc_interface4_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank4_core_initiator_length0_re = ((hdmi2usbsoc_csrbank4_sel & hdmi2usbsoc_interface4_bank_bus_we) & (hdmi2usbsoc_interface4_bank_bus_adr[4:0] == 5'd30));
assign hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage = hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage_full;
assign hdmi2usbsoc_csrbank4_core_underflow_enable0_w = hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage_full;
assign hdmi2usbsoc_csrbank4_core_underflow_counter3_w = hdmi2usbsoc_hdmi_out1_core_underflow_counter_status[31:24];
assign hdmi2usbsoc_csrbank4_core_underflow_counter2_w = hdmi2usbsoc_hdmi_out1_core_underflow_counter_status[23:16];
assign hdmi2usbsoc_csrbank4_core_underflow_counter1_w = hdmi2usbsoc_hdmi_out1_core_underflow_counter_status[15:8];
assign hdmi2usbsoc_csrbank4_core_underflow_counter0_w = hdmi2usbsoc_hdmi_out1_core_underflow_counter_status[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage = hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage_full;
assign hdmi2usbsoc_csrbank4_core_initiator_enable0_w = hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage_full;
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hres1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_hres0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_hscan1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_hscan0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vres1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_vres0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage_full[11:0];
assign hdmi2usbsoc_csrbank4_core_initiator_vscan1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage_full[11:8];
assign hdmi2usbsoc_csrbank4_core_initiator_vscan0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full[31:0];
assign hdmi2usbsoc_csrbank4_core_initiator_base3_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full[31:24];
assign hdmi2usbsoc_csrbank4_core_initiator_base2_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full[23:16];
assign hdmi2usbsoc_csrbank4_core_initiator_base1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full[15:8];
assign hdmi2usbsoc_csrbank4_core_initiator_base0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full[7:0];
assign hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full[31:0];
assign hdmi2usbsoc_csrbank4_core_initiator_length3_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full[31:24];
assign hdmi2usbsoc_csrbank4_core_initiator_length2_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full[23:16];
assign hdmi2usbsoc_csrbank4_core_initiator_length1_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full[15:8];
assign hdmi2usbsoc_csrbank4_core_initiator_length0_w = hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full[7:0];
assign hdmi2usbsoc_sram2_sel = (hdmi2usbsoc_interface2_sram_bus_adr[13:9] == 2'd3);

// synthesis translate_off
reg dummy_d_147;
// synthesis translate_on
always @(*) begin
	hdmi2usbsoc_interface2_sram_bus_dat_r <= 8'd0;
	if (hdmi2usbsoc_sram2_sel_r) begin
		hdmi2usbsoc_interface2_sram_bus_dat_r <= hdmi2usbsoc_sram2_dat_r;
	end
// synthesis translate_off
	dummy_d_147 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_sram2_adr = hdmi2usbsoc_interface2_sram_bus_adr[3:0];
assign hdmi2usbsoc_csrbank5_sel = (hdmi2usbsoc_interface5_bank_bus_adr[13:9] == 4'd12);
assign hdmi2usbsoc_csrbank5_dna_id7_r = hdmi2usbsoc_interface5_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank5_dna_id7_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 1'd0));
assign hdmi2usbsoc_csrbank5_dna_id6_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_dna_id6_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 1'd1));
assign hdmi2usbsoc_csrbank5_dna_id5_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_dna_id5_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 2'd2));
assign hdmi2usbsoc_csrbank5_dna_id4_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_dna_id4_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 2'd3));
assign hdmi2usbsoc_csrbank5_dna_id3_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_dna_id3_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 3'd4));
assign hdmi2usbsoc_csrbank5_dna_id2_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_dna_id2_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 3'd5));
assign hdmi2usbsoc_csrbank5_dna_id1_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_dna_id1_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 3'd6));
assign hdmi2usbsoc_csrbank5_dna_id0_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_dna_id0_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 3'd7));
assign hdmi2usbsoc_csrbank5_git_commit19_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit19_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd8));
assign hdmi2usbsoc_csrbank5_git_commit18_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit18_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd9));
assign hdmi2usbsoc_csrbank5_git_commit17_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit17_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd10));
assign hdmi2usbsoc_csrbank5_git_commit16_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit16_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd11));
assign hdmi2usbsoc_csrbank5_git_commit15_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit15_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd12));
assign hdmi2usbsoc_csrbank5_git_commit14_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit14_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd13));
assign hdmi2usbsoc_csrbank5_git_commit13_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit13_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd14));
assign hdmi2usbsoc_csrbank5_git_commit12_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit12_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 4'd15));
assign hdmi2usbsoc_csrbank5_git_commit11_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit11_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd16));
assign hdmi2usbsoc_csrbank5_git_commit10_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit10_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd17));
assign hdmi2usbsoc_csrbank5_git_commit9_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit9_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd18));
assign hdmi2usbsoc_csrbank5_git_commit8_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit8_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd19));
assign hdmi2usbsoc_csrbank5_git_commit7_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit7_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd20));
assign hdmi2usbsoc_csrbank5_git_commit6_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit6_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd21));
assign hdmi2usbsoc_csrbank5_git_commit5_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit5_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd22));
assign hdmi2usbsoc_csrbank5_git_commit4_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit4_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd23));
assign hdmi2usbsoc_csrbank5_git_commit3_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit3_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd24));
assign hdmi2usbsoc_csrbank5_git_commit2_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit2_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd25));
assign hdmi2usbsoc_csrbank5_git_commit1_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit1_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd26));
assign hdmi2usbsoc_csrbank5_git_commit0_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_git_commit0_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd27));
assign hdmi2usbsoc_csrbank5_platform_platform7_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform7_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd28));
assign hdmi2usbsoc_csrbank5_platform_platform6_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform6_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd29));
assign hdmi2usbsoc_csrbank5_platform_platform5_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform5_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd30));
assign hdmi2usbsoc_csrbank5_platform_platform4_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform4_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 5'd31));
assign hdmi2usbsoc_csrbank5_platform_platform3_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform3_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd32));
assign hdmi2usbsoc_csrbank5_platform_platform2_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform2_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd33));
assign hdmi2usbsoc_csrbank5_platform_platform1_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform1_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd34));
assign hdmi2usbsoc_csrbank5_platform_platform0_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform0_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd35));
assign hdmi2usbsoc_csrbank5_platform_target7_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target7_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd36));
assign hdmi2usbsoc_csrbank5_platform_target6_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target6_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd37));
assign hdmi2usbsoc_csrbank5_platform_target5_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target5_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd38));
assign hdmi2usbsoc_csrbank5_platform_target4_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target4_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd39));
assign hdmi2usbsoc_csrbank5_platform_target3_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target3_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd40));
assign hdmi2usbsoc_csrbank5_platform_target2_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target2_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd41));
assign hdmi2usbsoc_csrbank5_platform_target1_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target1_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd42));
assign hdmi2usbsoc_csrbank5_platform_target0_r = hdmi2usbsoc_interface5_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank5_platform_target0_re = ((hdmi2usbsoc_csrbank5_sel & hdmi2usbsoc_interface5_bank_bus_we) & (hdmi2usbsoc_interface5_bank_bus_adr[5:0] == 6'd43));
assign hdmi2usbsoc_csrbank5_dna_id7_w = hdmi2usbsoc_dna_status[56];
assign hdmi2usbsoc_csrbank5_dna_id6_w = hdmi2usbsoc_dna_status[55:48];
assign hdmi2usbsoc_csrbank5_dna_id5_w = hdmi2usbsoc_dna_status[47:40];
assign hdmi2usbsoc_csrbank5_dna_id4_w = hdmi2usbsoc_dna_status[39:32];
assign hdmi2usbsoc_csrbank5_dna_id3_w = hdmi2usbsoc_dna_status[31:24];
assign hdmi2usbsoc_csrbank5_dna_id2_w = hdmi2usbsoc_dna_status[23:16];
assign hdmi2usbsoc_csrbank5_dna_id1_w = hdmi2usbsoc_dna_status[15:8];
assign hdmi2usbsoc_csrbank5_dna_id0_w = hdmi2usbsoc_dna_status[7:0];
assign hdmi2usbsoc_csrbank5_git_commit19_w = hdmi2usbsoc_git_status[159:152];
assign hdmi2usbsoc_csrbank5_git_commit18_w = hdmi2usbsoc_git_status[151:144];
assign hdmi2usbsoc_csrbank5_git_commit17_w = hdmi2usbsoc_git_status[143:136];
assign hdmi2usbsoc_csrbank5_git_commit16_w = hdmi2usbsoc_git_status[135:128];
assign hdmi2usbsoc_csrbank5_git_commit15_w = hdmi2usbsoc_git_status[127:120];
assign hdmi2usbsoc_csrbank5_git_commit14_w = hdmi2usbsoc_git_status[119:112];
assign hdmi2usbsoc_csrbank5_git_commit13_w = hdmi2usbsoc_git_status[111:104];
assign hdmi2usbsoc_csrbank5_git_commit12_w = hdmi2usbsoc_git_status[103:96];
assign hdmi2usbsoc_csrbank5_git_commit11_w = hdmi2usbsoc_git_status[95:88];
assign hdmi2usbsoc_csrbank5_git_commit10_w = hdmi2usbsoc_git_status[87:80];
assign hdmi2usbsoc_csrbank5_git_commit9_w = hdmi2usbsoc_git_status[79:72];
assign hdmi2usbsoc_csrbank5_git_commit8_w = hdmi2usbsoc_git_status[71:64];
assign hdmi2usbsoc_csrbank5_git_commit7_w = hdmi2usbsoc_git_status[63:56];
assign hdmi2usbsoc_csrbank5_git_commit6_w = hdmi2usbsoc_git_status[55:48];
assign hdmi2usbsoc_csrbank5_git_commit5_w = hdmi2usbsoc_git_status[47:40];
assign hdmi2usbsoc_csrbank5_git_commit4_w = hdmi2usbsoc_git_status[39:32];
assign hdmi2usbsoc_csrbank5_git_commit3_w = hdmi2usbsoc_git_status[31:24];
assign hdmi2usbsoc_csrbank5_git_commit2_w = hdmi2usbsoc_git_status[23:16];
assign hdmi2usbsoc_csrbank5_git_commit1_w = hdmi2usbsoc_git_status[15:8];
assign hdmi2usbsoc_csrbank5_git_commit0_w = hdmi2usbsoc_git_status[7:0];
assign hdmi2usbsoc_csrbank5_platform_platform7_w = hdmi2usbsoc_platform_status[63:56];
assign hdmi2usbsoc_csrbank5_platform_platform6_w = hdmi2usbsoc_platform_status[55:48];
assign hdmi2usbsoc_csrbank5_platform_platform5_w = hdmi2usbsoc_platform_status[47:40];
assign hdmi2usbsoc_csrbank5_platform_platform4_w = hdmi2usbsoc_platform_status[39:32];
assign hdmi2usbsoc_csrbank5_platform_platform3_w = hdmi2usbsoc_platform_status[31:24];
assign hdmi2usbsoc_csrbank5_platform_platform2_w = hdmi2usbsoc_platform_status[23:16];
assign hdmi2usbsoc_csrbank5_platform_platform1_w = hdmi2usbsoc_platform_status[15:8];
assign hdmi2usbsoc_csrbank5_platform_platform0_w = hdmi2usbsoc_platform_status[7:0];
assign hdmi2usbsoc_csrbank5_platform_target7_w = hdmi2usbsoc_target_status[63:56];
assign hdmi2usbsoc_csrbank5_platform_target6_w = hdmi2usbsoc_target_status[55:48];
assign hdmi2usbsoc_csrbank5_platform_target5_w = hdmi2usbsoc_target_status[47:40];
assign hdmi2usbsoc_csrbank5_platform_target4_w = hdmi2usbsoc_target_status[39:32];
assign hdmi2usbsoc_csrbank5_platform_target3_w = hdmi2usbsoc_target_status[31:24];
assign hdmi2usbsoc_csrbank5_platform_target2_w = hdmi2usbsoc_target_status[23:16];
assign hdmi2usbsoc_csrbank5_platform_target1_w = hdmi2usbsoc_target_status[15:8];
assign hdmi2usbsoc_csrbank5_platform_target0_w = hdmi2usbsoc_target_status[7:0];
assign hdmi2usbsoc_csrbank6_sel = (hdmi2usbsoc_interface6_bank_bus_adr[13:9] == 4'd8);
assign hdmi2usbsoc_csrbank6_dfii_control0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank6_dfii_control0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 1'd0));
assign hdmi2usbsoc_csrbank6_dfii_pi0_command0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_command0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 1'd1));
assign hdmi2usbsoc_sdram_phaseinjector0_command_issue_r = hdmi2usbsoc_interface6_bank_bus_dat_w[0];
assign hdmi2usbsoc_sdram_phaseinjector0_command_issue_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 2'd2));
assign hdmi2usbsoc_csrbank6_dfii_pi0_address1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[4:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_address1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 2'd3));
assign hdmi2usbsoc_csrbank6_dfii_pi0_address0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_address0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 3'd4));
assign hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 3'd5));
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 3'd6));
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 3'd7));
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd8));
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd9));
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata3_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata3_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd10));
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata2_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata2_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd11));
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd12));
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd13));
assign hdmi2usbsoc_csrbank6_dfii_pi1_command0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[5:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_command0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd14));
assign hdmi2usbsoc_sdram_phaseinjector1_command_issue_r = hdmi2usbsoc_interface6_bank_bus_dat_w[0];
assign hdmi2usbsoc_sdram_phaseinjector1_command_issue_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 4'd15));
assign hdmi2usbsoc_csrbank6_dfii_pi1_address1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[4:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_address1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd16));
assign hdmi2usbsoc_csrbank6_dfii_pi1_address0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_address0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd17));
assign hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[2:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd18));
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd19));
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd20));
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd21));
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd22));
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata3_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata3_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd23));
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata2_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata2_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd24));
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd25));
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd26));
assign hdmi2usbsoc_sdram_bandwidth_update_r = hdmi2usbsoc_interface6_bank_bus_dat_w[0];
assign hdmi2usbsoc_sdram_bandwidth_update_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd27));
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads2_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads2_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd28));
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd29));
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd30));
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites2_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites2_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 5'd31));
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites1_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites1_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 6'd32));
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites0_r = hdmi2usbsoc_interface6_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites0_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 6'd33));
assign hdmi2usbsoc_csrbank6_controller_bandwidth_data_width_r = hdmi2usbsoc_interface6_bank_bus_dat_w[6:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_data_width_re = ((hdmi2usbsoc_csrbank6_sel & hdmi2usbsoc_interface6_bank_bus_we) & (hdmi2usbsoc_interface6_bank_bus_adr[5:0] == 6'd34));
assign hdmi2usbsoc_sdram_storage = hdmi2usbsoc_sdram_storage_full[3:0];
assign hdmi2usbsoc_csrbank6_dfii_control0_w = hdmi2usbsoc_sdram_storage_full[3:0];
assign hdmi2usbsoc_sdram_phaseinjector0_command_storage = hdmi2usbsoc_sdram_phaseinjector0_command_storage_full[5:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_command0_w = hdmi2usbsoc_sdram_phaseinjector0_command_storage_full[5:0];
assign hdmi2usbsoc_sdram_phaseinjector0_address_storage = hdmi2usbsoc_sdram_phaseinjector0_address_storage_full[12:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_address1_w = hdmi2usbsoc_sdram_phaseinjector0_address_storage_full[12:8];
assign hdmi2usbsoc_csrbank6_dfii_pi0_address0_w = hdmi2usbsoc_sdram_phaseinjector0_address_storage_full[7:0];
assign hdmi2usbsoc_sdram_phaseinjector0_baddress_storage = hdmi2usbsoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_w = hdmi2usbsoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage = hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[31:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_w = hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[31:24];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_w = hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[23:16];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_w = hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[15:8];
assign hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_w = hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata3_w = hdmi2usbsoc_sdram_phaseinjector0_status[31:24];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata2_w = hdmi2usbsoc_sdram_phaseinjector0_status[23:16];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata1_w = hdmi2usbsoc_sdram_phaseinjector0_status[15:8];
assign hdmi2usbsoc_csrbank6_dfii_pi0_rddata0_w = hdmi2usbsoc_sdram_phaseinjector0_status[7:0];
assign hdmi2usbsoc_sdram_phaseinjector1_command_storage = hdmi2usbsoc_sdram_phaseinjector1_command_storage_full[5:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_command0_w = hdmi2usbsoc_sdram_phaseinjector1_command_storage_full[5:0];
assign hdmi2usbsoc_sdram_phaseinjector1_address_storage = hdmi2usbsoc_sdram_phaseinjector1_address_storage_full[12:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_address1_w = hdmi2usbsoc_sdram_phaseinjector1_address_storage_full[12:8];
assign hdmi2usbsoc_csrbank6_dfii_pi1_address0_w = hdmi2usbsoc_sdram_phaseinjector1_address_storage_full[7:0];
assign hdmi2usbsoc_sdram_phaseinjector1_baddress_storage = hdmi2usbsoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_w = hdmi2usbsoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage = hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[31:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_w = hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[31:24];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_w = hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[23:16];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_w = hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[15:8];
assign hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_w = hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[7:0];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata3_w = hdmi2usbsoc_sdram_phaseinjector1_status[31:24];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata2_w = hdmi2usbsoc_sdram_phaseinjector1_status[23:16];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata1_w = hdmi2usbsoc_sdram_phaseinjector1_status[15:8];
assign hdmi2usbsoc_csrbank6_dfii_pi1_rddata0_w = hdmi2usbsoc_sdram_phaseinjector1_status[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads2_w = hdmi2usbsoc_sdram_bandwidth_nreads_status[23:16];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads1_w = hdmi2usbsoc_sdram_bandwidth_nreads_status[15:8];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nreads0_w = hdmi2usbsoc_sdram_bandwidth_nreads_status[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites2_w = hdmi2usbsoc_sdram_bandwidth_nwrites_status[23:16];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites1_w = hdmi2usbsoc_sdram_bandwidth_nwrites_status[15:8];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites0_w = hdmi2usbsoc_sdram_bandwidth_nwrites_status[7:0];
assign hdmi2usbsoc_csrbank6_controller_bandwidth_data_width_w = hdmi2usbsoc_sdram_bandwidth_data_width_status[6:0];
assign hdmi2usbsoc_csrbank7_sel = (hdmi2usbsoc_interface7_bank_bus_adr[13:9] == 4'd10);
assign hdmi2usbsoc_csrbank7_bitbang0_r = hdmi2usbsoc_interface7_bank_bus_dat_w[3:0];
assign hdmi2usbsoc_csrbank7_bitbang0_re = ((hdmi2usbsoc_csrbank7_sel & hdmi2usbsoc_interface7_bank_bus_we) & (hdmi2usbsoc_interface7_bank_bus_adr[1:0] == 1'd0));
assign hdmi2usbsoc_csrbank7_miso_r = hdmi2usbsoc_interface7_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank7_miso_re = ((hdmi2usbsoc_csrbank7_sel & hdmi2usbsoc_interface7_bank_bus_we) & (hdmi2usbsoc_interface7_bank_bus_adr[1:0] == 1'd1));
assign hdmi2usbsoc_csrbank7_bitbang_en0_r = hdmi2usbsoc_interface7_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank7_bitbang_en0_re = ((hdmi2usbsoc_csrbank7_sel & hdmi2usbsoc_interface7_bank_bus_we) & (hdmi2usbsoc_interface7_bank_bus_adr[1:0] == 2'd2));
assign hdmi2usbsoc_bitbang_storage = hdmi2usbsoc_bitbang_storage_full[3:0];
assign hdmi2usbsoc_csrbank7_bitbang0_w = hdmi2usbsoc_bitbang_storage_full[3:0];
assign hdmi2usbsoc_csrbank7_miso_w = hdmi2usbsoc_status;
assign hdmi2usbsoc_bitbang_en_storage = hdmi2usbsoc_bitbang_en_storage_full;
assign hdmi2usbsoc_csrbank7_bitbang_en0_w = hdmi2usbsoc_bitbang_en_storage_full;
assign hdmi2usbsoc_csrbank8_sel = (hdmi2usbsoc_interface8_bank_bus_adr[13:9] == 3'd4);
assign hdmi2usbsoc_csrbank8_load3_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_load3_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 1'd0));
assign hdmi2usbsoc_csrbank8_load2_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_load2_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 1'd1));
assign hdmi2usbsoc_csrbank8_load1_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_load1_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 2'd2));
assign hdmi2usbsoc_csrbank8_load0_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_load0_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 2'd3));
assign hdmi2usbsoc_csrbank8_reload3_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_reload3_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 3'd4));
assign hdmi2usbsoc_csrbank8_reload2_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_reload2_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 3'd5));
assign hdmi2usbsoc_csrbank8_reload1_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_reload1_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 3'd6));
assign hdmi2usbsoc_csrbank8_reload0_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_reload0_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 3'd7));
assign hdmi2usbsoc_csrbank8_en0_r = hdmi2usbsoc_interface8_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank8_en0_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd8));
assign hdmi2usbsoc_hdmi2usbsoc_timer0_update_value_r = hdmi2usbsoc_interface8_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi2usbsoc_timer0_update_value_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd9));
assign hdmi2usbsoc_csrbank8_value3_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_value3_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd10));
assign hdmi2usbsoc_csrbank8_value2_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_value2_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd11));
assign hdmi2usbsoc_csrbank8_value1_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_value1_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd12));
assign hdmi2usbsoc_csrbank8_value0_r = hdmi2usbsoc_interface8_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank8_value0_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd13));
assign hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_status_r = hdmi2usbsoc_interface8_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_status_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd14));
assign hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_r = hdmi2usbsoc_interface8_bank_bus_dat_w[0];
assign hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 4'd15));
assign hdmi2usbsoc_csrbank8_ev_enable0_r = hdmi2usbsoc_interface8_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank8_ev_enable0_re = ((hdmi2usbsoc_csrbank8_sel & hdmi2usbsoc_interface8_bank_bus_we) & (hdmi2usbsoc_interface8_bank_bus_adr[4:0] == 5'd16));
assign hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage = hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[31:0];
assign hdmi2usbsoc_csrbank8_load3_w = hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[31:24];
assign hdmi2usbsoc_csrbank8_load2_w = hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[23:16];
assign hdmi2usbsoc_csrbank8_load1_w = hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[15:8];
assign hdmi2usbsoc_csrbank8_load0_w = hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[7:0];
assign hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage = hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[31:0];
assign hdmi2usbsoc_csrbank8_reload3_w = hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[31:24];
assign hdmi2usbsoc_csrbank8_reload2_w = hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[23:16];
assign hdmi2usbsoc_csrbank8_reload1_w = hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[15:8];
assign hdmi2usbsoc_csrbank8_reload0_w = hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[7:0];
assign hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage = hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage_full;
assign hdmi2usbsoc_csrbank8_en0_w = hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage_full;
assign hdmi2usbsoc_csrbank8_value3_w = hdmi2usbsoc_hdmi2usbsoc_timer0_value_status[31:24];
assign hdmi2usbsoc_csrbank8_value2_w = hdmi2usbsoc_hdmi2usbsoc_timer0_value_status[23:16];
assign hdmi2usbsoc_csrbank8_value1_w = hdmi2usbsoc_hdmi2usbsoc_timer0_value_status[15:8];
assign hdmi2usbsoc_csrbank8_value0_w = hdmi2usbsoc_hdmi2usbsoc_timer0_value_status[7:0];
assign hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage = hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage_full;
assign hdmi2usbsoc_csrbank8_ev_enable0_w = hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage_full;
assign hdmi2usbsoc_csrbank9_sel = (hdmi2usbsoc_interface9_bank_bus_adr[13:9] == 2'd2);
assign hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_r = hdmi2usbsoc_interface9_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_re = ((hdmi2usbsoc_csrbank9_sel & hdmi2usbsoc_interface9_bank_bus_we) & (hdmi2usbsoc_interface9_bank_bus_adr[2:0] == 1'd0));
assign hdmi2usbsoc_csrbank9_txfull_r = hdmi2usbsoc_interface9_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank9_txfull_re = ((hdmi2usbsoc_csrbank9_sel & hdmi2usbsoc_interface9_bank_bus_we) & (hdmi2usbsoc_interface9_bank_bus_adr[2:0] == 1'd1));
assign hdmi2usbsoc_csrbank9_rxempty_r = hdmi2usbsoc_interface9_bank_bus_dat_w[0];
assign hdmi2usbsoc_csrbank9_rxempty_re = ((hdmi2usbsoc_csrbank9_sel & hdmi2usbsoc_interface9_bank_bus_we) & (hdmi2usbsoc_interface9_bank_bus_adr[2:0] == 2'd2));
assign hdmi2usbsoc_hdmi2usbsoc_uart_status_r = hdmi2usbsoc_interface9_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_hdmi2usbsoc_uart_status_re = ((hdmi2usbsoc_csrbank9_sel & hdmi2usbsoc_interface9_bank_bus_we) & (hdmi2usbsoc_interface9_bank_bus_adr[2:0] == 2'd3));
assign hdmi2usbsoc_hdmi2usbsoc_uart_pending_r = hdmi2usbsoc_interface9_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_hdmi2usbsoc_uart_pending_re = ((hdmi2usbsoc_csrbank9_sel & hdmi2usbsoc_interface9_bank_bus_we) & (hdmi2usbsoc_interface9_bank_bus_adr[2:0] == 3'd4));
assign hdmi2usbsoc_csrbank9_ev_enable0_r = hdmi2usbsoc_interface9_bank_bus_dat_w[1:0];
assign hdmi2usbsoc_csrbank9_ev_enable0_re = ((hdmi2usbsoc_csrbank9_sel & hdmi2usbsoc_interface9_bank_bus_we) & (hdmi2usbsoc_interface9_bank_bus_adr[2:0] == 3'd5));
assign hdmi2usbsoc_csrbank9_txfull_w = hdmi2usbsoc_hdmi2usbsoc_uart_txfull_status;
assign hdmi2usbsoc_csrbank9_rxempty_w = hdmi2usbsoc_hdmi2usbsoc_uart_rxempty_status;
assign hdmi2usbsoc_hdmi2usbsoc_uart_storage = hdmi2usbsoc_hdmi2usbsoc_uart_storage_full[1:0];
assign hdmi2usbsoc_csrbank9_ev_enable0_w = hdmi2usbsoc_hdmi2usbsoc_uart_storage_full[1:0];
assign hdmi2usbsoc_csrbank10_sel = (hdmi2usbsoc_interface10_bank_bus_adr[13:9] == 1'd1);
assign hdmi2usbsoc_csrbank10_tuning_word3_r = hdmi2usbsoc_interface10_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank10_tuning_word3_re = ((hdmi2usbsoc_csrbank10_sel & hdmi2usbsoc_interface10_bank_bus_we) & (hdmi2usbsoc_interface10_bank_bus_adr[1:0] == 1'd0));
assign hdmi2usbsoc_csrbank10_tuning_word2_r = hdmi2usbsoc_interface10_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank10_tuning_word2_re = ((hdmi2usbsoc_csrbank10_sel & hdmi2usbsoc_interface10_bank_bus_we) & (hdmi2usbsoc_interface10_bank_bus_adr[1:0] == 1'd1));
assign hdmi2usbsoc_csrbank10_tuning_word1_r = hdmi2usbsoc_interface10_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank10_tuning_word1_re = ((hdmi2usbsoc_csrbank10_sel & hdmi2usbsoc_interface10_bank_bus_we) & (hdmi2usbsoc_interface10_bank_bus_adr[1:0] == 2'd2));
assign hdmi2usbsoc_csrbank10_tuning_word0_r = hdmi2usbsoc_interface10_bank_bus_dat_w[7:0];
assign hdmi2usbsoc_csrbank10_tuning_word0_re = ((hdmi2usbsoc_csrbank10_sel & hdmi2usbsoc_interface10_bank_bus_we) & (hdmi2usbsoc_interface10_bank_bus_adr[1:0] == 2'd3));
assign hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage = hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[31:0];
assign hdmi2usbsoc_csrbank10_tuning_word3_w = hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[31:24];
assign hdmi2usbsoc_csrbank10_tuning_word2_w = hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[23:16];
assign hdmi2usbsoc_csrbank10_tuning_word1_w = hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[15:8];
assign hdmi2usbsoc_csrbank10_tuning_word0_w = hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[7:0];
assign hdmi2usbsoc_interface0_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface1_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface2_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface3_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface4_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface5_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface6_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface7_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface8_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface9_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface10_bank_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface0_sram_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface1_sram_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface2_sram_bus_adr = hdmi2usbsoc_hdmi2usbsoc_interface_adr;
assign hdmi2usbsoc_interface0_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface1_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface2_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface3_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface4_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface5_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface6_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface7_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface8_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface9_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface10_bank_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface0_sram_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface1_sram_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface2_sram_bus_we = hdmi2usbsoc_hdmi2usbsoc_interface_we;
assign hdmi2usbsoc_interface0_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface1_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface2_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface3_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface4_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface5_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface6_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface7_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface8_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface9_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface10_bank_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface0_sram_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface1_sram_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_interface2_sram_bus_dat_w = hdmi2usbsoc_hdmi2usbsoc_interface_dat_w;
assign hdmi2usbsoc_hdmi2usbsoc_interface_dat_r = (((((((((((((hdmi2usbsoc_interface0_bank_bus_dat_r | hdmi2usbsoc_interface1_bank_bus_dat_r) | hdmi2usbsoc_interface2_bank_bus_dat_r) | hdmi2usbsoc_interface3_bank_bus_dat_r) | hdmi2usbsoc_interface4_bank_bus_dat_r) | hdmi2usbsoc_interface5_bank_bus_dat_r) | hdmi2usbsoc_interface6_bank_bus_dat_r) | hdmi2usbsoc_interface7_bank_bus_dat_r) | hdmi2usbsoc_interface8_bank_bus_dat_r) | hdmi2usbsoc_interface9_bank_bus_dat_r) | hdmi2usbsoc_interface10_bank_bus_dat_r) | hdmi2usbsoc_interface0_sram_bus_dat_r) | hdmi2usbsoc_interface1_sram_bus_dat_r) | hdmi2usbsoc_interface2_sram_bus_dat_r);
assign slice_proxy0 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy1 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy2 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy3 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy4 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy5 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy6 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy7 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy8 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy9 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy10 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy11 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy12 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy13 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy14 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy15 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy16 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy17 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy18 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy19 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy20 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy21 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy22 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy23 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy24 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy25 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy26 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy27 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy28 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy29 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy30 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy31 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy32 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy33 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy34 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy35 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy36 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy37 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy38 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy39 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy40 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy41 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy42 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy43 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy44 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy45 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy46 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy47 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy48 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy49 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy50 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy51 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy52 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy53 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy54 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy55 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy56 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy57 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy58 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy59 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy60 = hdmi2usbsoc_ddrphy_record2_wrdata[31:16];
assign slice_proxy61 = hdmi2usbsoc_ddrphy_record2_wrdata[15:0];
assign slice_proxy62 = hdmi2usbsoc_ddrphy_record3_wrdata[31:16];
assign slice_proxy63 = hdmi2usbsoc_ddrphy_record3_wrdata[15:0];
assign slice_proxy64 = hdmi2usbsoc_ddrphy_record2_wrdata_mask[3:2];
assign slice_proxy65 = hdmi2usbsoc_ddrphy_record2_wrdata_mask[1:0];
assign slice_proxy66 = hdmi2usbsoc_ddrphy_record3_wrdata_mask[3:2];
assign slice_proxy67 = hdmi2usbsoc_ddrphy_record3_wrdata_mask[1:0];
assign slice_proxy68 = hdmi2usbsoc_ddrphy_record2_wrdata_mask[3:2];
assign slice_proxy69 = hdmi2usbsoc_ddrphy_record2_wrdata_mask[1:0];
assign slice_proxy70 = hdmi2usbsoc_ddrphy_record3_wrdata_mask[3:2];
assign slice_proxy71 = hdmi2usbsoc_ddrphy_record3_wrdata_mask[1:0];

// synthesis translate_off
reg dummy_d_148;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed0 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[0];
		end
		1'd1: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[1];
		end
		2'd2: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[2];
		end
		2'd3: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[3];
		end
		3'd4: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[4];
		end
		3'd5: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[5];
		end
		3'd6: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[6];
		end
		default: begin
			comb_rhs_array_muxed0 <= hdmi2usbsoc_sdram_choose_cmd_valids[7];
		end
	endcase
// synthesis translate_off
	dummy_d_148 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_149;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed1 <= 13'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			comb_rhs_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
// synthesis translate_off
	dummy_d_149 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_150;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed2 <= 3'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			comb_rhs_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
// synthesis translate_off
	dummy_d_150 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_151;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed3 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			comb_rhs_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
// synthesis translate_off
	dummy_d_151 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_152;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed4 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			comb_rhs_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
// synthesis translate_off
	dummy_d_152 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_153;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed5 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			comb_rhs_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
// synthesis translate_off
	dummy_d_153 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_154;
// synthesis translate_on
always @(*) begin
	comb_t_array_muxed0 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			comb_t_array_muxed0 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
// synthesis translate_off
	dummy_d_154 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_155;
// synthesis translate_on
always @(*) begin
	comb_t_array_muxed1 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			comb_t_array_muxed1 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
// synthesis translate_off
	dummy_d_155 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_156;
// synthesis translate_on
always @(*) begin
	comb_t_array_muxed2 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_cmd_grant)
		1'd0: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			comb_t_array_muxed2 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_156 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_157;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed6 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[0];
		end
		1'd1: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[1];
		end
		2'd2: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[2];
		end
		2'd3: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[3];
		end
		3'd4: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[4];
		end
		3'd5: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[5];
		end
		3'd6: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[6];
		end
		default: begin
			comb_rhs_array_muxed6 <= hdmi2usbsoc_sdram_choose_req_valids[7];
		end
	endcase
// synthesis translate_off
	dummy_d_157 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_158;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed7 <= 13'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			comb_rhs_array_muxed7 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
// synthesis translate_off
	dummy_d_158 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_159;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed8 <= 3'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			comb_rhs_array_muxed8 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
// synthesis translate_off
	dummy_d_159 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_160;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed9 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			comb_rhs_array_muxed9 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
// synthesis translate_off
	dummy_d_160 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_161;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed10 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			comb_rhs_array_muxed10 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
// synthesis translate_off
	dummy_d_161 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_162;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed11 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			comb_rhs_array_muxed11 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
// synthesis translate_off
	dummy_d_162 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_163;
// synthesis translate_on
always @(*) begin
	comb_t_array_muxed3 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			comb_t_array_muxed3 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
// synthesis translate_off
	dummy_d_163 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_164;
// synthesis translate_on
always @(*) begin
	comb_t_array_muxed4 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			comb_t_array_muxed4 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
// synthesis translate_off
	dummy_d_164 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_165;
// synthesis translate_on
always @(*) begin
	comb_t_array_muxed5 <= 1'd0;
	case (hdmi2usbsoc_sdram_choose_req_grant)
		1'd0: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			comb_t_array_muxed5 <= hdmi2usbsoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_165 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_166;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed12 <= 21'd0;
	case (controllerinjector_roundrobin0_grant)
		1'd0: begin
			comb_rhs_array_muxed12 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed12 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed12 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed12 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed12 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed12 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_166 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_167;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed13 <= 1'd0;
	case (controllerinjector_roundrobin0_grant)
		1'd0: begin
			comb_rhs_array_muxed13 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed13 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed13 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed13 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed13 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed13 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_167 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_168;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed14 <= 1'd0;
	case (controllerinjector_roundrobin0_grant)
		1'd0: begin
			comb_rhs_array_muxed14 <= (((controllerinjector_cba0 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed14 <= (((controllerinjector_cba1 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed14 <= (((controllerinjector_cba2 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed14 <= (((controllerinjector_cba3 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed14 <= (((controllerinjector_cba4 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed14 <= (((controllerinjector_cba5 == 1'd0) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_168 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_169;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed15 <= 21'd0;
	case (controllerinjector_roundrobin1_grant)
		1'd0: begin
			comb_rhs_array_muxed15 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed15 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed15 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed15 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed15 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed15 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_169 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_170;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed16 <= 1'd0;
	case (controllerinjector_roundrobin1_grant)
		1'd0: begin
			comb_rhs_array_muxed16 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed16 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed16 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed16 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed16 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed16 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_170 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_171;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed17 <= 1'd0;
	case (controllerinjector_roundrobin1_grant)
		1'd0: begin
			comb_rhs_array_muxed17 <= (((controllerinjector_cba0 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed17 <= (((controllerinjector_cba1 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed17 <= (((controllerinjector_cba2 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed17 <= (((controllerinjector_cba3 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed17 <= (((controllerinjector_cba4 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed17 <= (((controllerinjector_cba5 == 1'd1) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_171 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_172;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed18 <= 21'd0;
	case (controllerinjector_roundrobin2_grant)
		1'd0: begin
			comb_rhs_array_muxed18 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed18 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed18 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed18 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed18 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed18 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_172 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_173;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed19 <= 1'd0;
	case (controllerinjector_roundrobin2_grant)
		1'd0: begin
			comb_rhs_array_muxed19 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed19 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed19 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed19 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed19 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed19 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_173 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_174;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed20 <= 1'd0;
	case (controllerinjector_roundrobin2_grant)
		1'd0: begin
			comb_rhs_array_muxed20 <= (((controllerinjector_cba0 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed20 <= (((controllerinjector_cba1 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed20 <= (((controllerinjector_cba2 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed20 <= (((controllerinjector_cba3 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed20 <= (((controllerinjector_cba4 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed20 <= (((controllerinjector_cba5 == 2'd2) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_174 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_175;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed21 <= 21'd0;
	case (controllerinjector_roundrobin3_grant)
		1'd0: begin
			comb_rhs_array_muxed21 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed21 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed21 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed21 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed21 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed21 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_175 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_176;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed22 <= 1'd0;
	case (controllerinjector_roundrobin3_grant)
		1'd0: begin
			comb_rhs_array_muxed22 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed22 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed22 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed22 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed22 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed22 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_176 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_177;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed23 <= 1'd0;
	case (controllerinjector_roundrobin3_grant)
		1'd0: begin
			comb_rhs_array_muxed23 <= (((controllerinjector_cba0 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed23 <= (((controllerinjector_cba1 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed23 <= (((controllerinjector_cba2 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed23 <= (((controllerinjector_cba3 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed23 <= (((controllerinjector_cba4 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed23 <= (((controllerinjector_cba5 == 2'd3) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_177 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_178;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed24 <= 21'd0;
	case (controllerinjector_roundrobin4_grant)
		1'd0: begin
			comb_rhs_array_muxed24 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed24 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed24 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed24 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed24 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed24 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_178 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_179;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed25 <= 1'd0;
	case (controllerinjector_roundrobin4_grant)
		1'd0: begin
			comb_rhs_array_muxed25 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed25 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed25 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed25 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed25 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed25 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_179 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_180;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed26 <= 1'd0;
	case (controllerinjector_roundrobin4_grant)
		1'd0: begin
			comb_rhs_array_muxed26 <= (((controllerinjector_cba0 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed26 <= (((controllerinjector_cba1 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed26 <= (((controllerinjector_cba2 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed26 <= (((controllerinjector_cba3 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed26 <= (((controllerinjector_cba4 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed26 <= (((controllerinjector_cba5 == 3'd4) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_180 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_181;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed27 <= 21'd0;
	case (controllerinjector_roundrobin5_grant)
		1'd0: begin
			comb_rhs_array_muxed27 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed27 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed27 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed27 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed27 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed27 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_181 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_182;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed28 <= 1'd0;
	case (controllerinjector_roundrobin5_grant)
		1'd0: begin
			comb_rhs_array_muxed28 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed28 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed28 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed28 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed28 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed28 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_182 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_183;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed29 <= 1'd0;
	case (controllerinjector_roundrobin5_grant)
		1'd0: begin
			comb_rhs_array_muxed29 <= (((controllerinjector_cba0 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed29 <= (((controllerinjector_cba1 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed29 <= (((controllerinjector_cba2 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed29 <= (((controllerinjector_cba3 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed29 <= (((controllerinjector_cba4 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed29 <= (((controllerinjector_cba5 == 3'd5) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_183 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_184;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed30 <= 21'd0;
	case (controllerinjector_roundrobin6_grant)
		1'd0: begin
			comb_rhs_array_muxed30 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed30 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed30 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed30 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed30 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed30 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_184 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_185;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed31 <= 1'd0;
	case (controllerinjector_roundrobin6_grant)
		1'd0: begin
			comb_rhs_array_muxed31 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed31 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed31 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed31 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed31 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed31 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_185 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_186;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed32 <= 1'd0;
	case (controllerinjector_roundrobin6_grant)
		1'd0: begin
			comb_rhs_array_muxed32 <= (((controllerinjector_cba0 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed32 <= (((controllerinjector_cba1 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed32 <= (((controllerinjector_cba2 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed32 <= (((controllerinjector_cba3 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed32 <= (((controllerinjector_cba4 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed32 <= (((controllerinjector_cba5 == 3'd6) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank7_lock & (controllerinjector_roundrobin7_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_186 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_187;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed33 <= 21'd0;
	case (controllerinjector_roundrobin7_grant)
		1'd0: begin
			comb_rhs_array_muxed33 <= controllerinjector_rca0;
		end
		1'd1: begin
			comb_rhs_array_muxed33 <= controllerinjector_rca1;
		end
		2'd2: begin
			comb_rhs_array_muxed33 <= controllerinjector_rca2;
		end
		2'd3: begin
			comb_rhs_array_muxed33 <= controllerinjector_rca3;
		end
		3'd4: begin
			comb_rhs_array_muxed33 <= controllerinjector_rca4;
		end
		default: begin
			comb_rhs_array_muxed33 <= controllerinjector_rca5;
		end
	endcase
// synthesis translate_off
	dummy_d_187 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_188;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed34 <= 1'd0;
	case (controllerinjector_roundrobin7_grant)
		1'd0: begin
			comb_rhs_array_muxed34 <= hdmi2usbsoc_port_cmd_payload_we;
		end
		1'd1: begin
			comb_rhs_array_muxed34 <= hdmi2usbsoc_litedramport0_cmd_payload_we0;
		end
		2'd2: begin
			comb_rhs_array_muxed34 <= hdmi2usbsoc_litedramport1_cmd_payload_we0;
		end
		2'd3: begin
			comb_rhs_array_muxed34 <= hdmi2usbsoc_litedramport2_cmd_payload_we0;
		end
		3'd4: begin
			comb_rhs_array_muxed34 <= hdmi2usbsoc_litedramport3_cmd_payload_we0;
		end
		default: begin
			comb_rhs_array_muxed34 <= encoder_port_port_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_188 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_189;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed35 <= 1'd0;
	case (controllerinjector_roundrobin7_grant)
		1'd0: begin
			comb_rhs_array_muxed35 <= (((controllerinjector_cba0 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd0))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd0))))) & hdmi2usbsoc_port_cmd_valid);
		end
		1'd1: begin
			comb_rhs_array_muxed35 <= (((controllerinjector_cba1 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 1'd1))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 1'd1))))) & hdmi2usbsoc_litedramport0_cmd_valid0);
		end
		2'd2: begin
			comb_rhs_array_muxed35 <= (((controllerinjector_cba2 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd2))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd2))))) & hdmi2usbsoc_litedramport1_cmd_valid0);
		end
		2'd3: begin
			comb_rhs_array_muxed35 <= (((controllerinjector_cba3 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 2'd3))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 2'd3))))) & hdmi2usbsoc_litedramport2_cmd_valid0);
		end
		3'd4: begin
			comb_rhs_array_muxed35 <= (((controllerinjector_cba4 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd4))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd4))))) & hdmi2usbsoc_litedramport3_cmd_valid0);
		end
		default: begin
			comb_rhs_array_muxed35 <= (((controllerinjector_cba5 == 3'd7) & (~(((((((1'd0 | (hdmi2usbsoc_sdram_interface_bank0_lock & (controllerinjector_roundrobin0_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank1_lock & (controllerinjector_roundrobin1_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank2_lock & (controllerinjector_roundrobin2_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank3_lock & (controllerinjector_roundrobin3_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank4_lock & (controllerinjector_roundrobin4_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank5_lock & (controllerinjector_roundrobin5_grant == 3'd5))) | (hdmi2usbsoc_sdram_interface_bank6_lock & (controllerinjector_roundrobin6_grant == 3'd5))))) & encoder_port_port_cmd_valid);
		end
	endcase
// synthesis translate_off
	dummy_d_189 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_190;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed36 <= 24'd0;
	case (hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot)
		1'd0: begin
			comb_rhs_array_muxed36 <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address;
		end
		default: begin
			comb_rhs_array_muxed36 <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address;
		end
	endcase
// synthesis translate_off
	dummy_d_190 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_191;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed37 <= 1'd0;
	case (hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot)
		1'd0: begin
			comb_rhs_array_muxed37 <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_valid;
		end
		default: begin
			comb_rhs_array_muxed37 <= hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_valid;
		end
	endcase
// synthesis translate_off
	dummy_d_191 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_192;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed38 <= 24'd0;
	case (hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot)
		1'd0: begin
			comb_rhs_array_muxed38 <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address;
		end
		default: begin
			comb_rhs_array_muxed38 <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address;
		end
	endcase
// synthesis translate_off
	dummy_d_192 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_193;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed39 <= 1'd0;
	case (hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot)
		1'd0: begin
			comb_rhs_array_muxed39 <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_valid;
		end
		default: begin
			comb_rhs_array_muxed39 <= hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_valid;
		end
	endcase
// synthesis translate_off
	dummy_d_193 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_194;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed40 <= 30'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed40 <= hdmi2usbsoc_interface1_wb_sdram_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_194 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_195;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed41 <= 32'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed41 <= hdmi2usbsoc_interface1_wb_sdram_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_195 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_196;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed42 <= 4'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed42 <= hdmi2usbsoc_interface1_wb_sdram_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_196 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_197;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed43 <= 1'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed43 <= hdmi2usbsoc_interface1_wb_sdram_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_197 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_198;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed44 <= 1'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed44 <= hdmi2usbsoc_interface1_wb_sdram_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_198 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_199;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed45 <= 1'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed45 <= hdmi2usbsoc_interface1_wb_sdram_we;
		end
	endcase
// synthesis translate_off
	dummy_d_199 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_200;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed46 <= 3'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed46 <= hdmi2usbsoc_interface1_wb_sdram_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_200 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_201;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed47 <= 2'd0;
	case (wb_sdram_con_grant)
		default: begin
			comb_rhs_array_muxed47 <= hdmi2usbsoc_interface1_wb_sdram_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_201 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_202;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed48 <= 30'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed48 <= hdmi2usbsoc_hdmi2usbsoc_ibus_adr;
		end
		default: begin
			comb_rhs_array_muxed48 <= hdmi2usbsoc_hdmi2usbsoc_dbus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_202 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_203;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed49 <= 32'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed49 <= hdmi2usbsoc_hdmi2usbsoc_ibus_dat_w;
		end
		default: begin
			comb_rhs_array_muxed49 <= hdmi2usbsoc_hdmi2usbsoc_dbus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_203 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_204;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed50 <= 4'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed50 <= hdmi2usbsoc_hdmi2usbsoc_ibus_sel;
		end
		default: begin
			comb_rhs_array_muxed50 <= hdmi2usbsoc_hdmi2usbsoc_dbus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_204 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_205;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed51 <= 1'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed51 <= hdmi2usbsoc_hdmi2usbsoc_ibus_cyc;
		end
		default: begin
			comb_rhs_array_muxed51 <= hdmi2usbsoc_hdmi2usbsoc_dbus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_205 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_206;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed52 <= 1'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed52 <= hdmi2usbsoc_hdmi2usbsoc_ibus_stb;
		end
		default: begin
			comb_rhs_array_muxed52 <= hdmi2usbsoc_hdmi2usbsoc_dbus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_206 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_207;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed53 <= 1'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed53 <= hdmi2usbsoc_hdmi2usbsoc_ibus_we;
		end
		default: begin
			comb_rhs_array_muxed53 <= hdmi2usbsoc_hdmi2usbsoc_dbus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_207 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_208;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed54 <= 3'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed54 <= hdmi2usbsoc_hdmi2usbsoc_ibus_cti;
		end
		default: begin
			comb_rhs_array_muxed54 <= hdmi2usbsoc_hdmi2usbsoc_dbus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_208 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_209;
// synthesis translate_on
always @(*) begin
	comb_rhs_array_muxed55 <= 2'd0;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			comb_rhs_array_muxed55 <= hdmi2usbsoc_hdmi2usbsoc_ibus_bte;
		end
		default: begin
			comb_rhs_array_muxed55 <= hdmi2usbsoc_hdmi2usbsoc_dbus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_209 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_210;
// synthesis translate_on
always @(*) begin
	sync_f_array_muxed0 <= 10'd0;
	case (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c2)
		1'd0: begin
			sync_f_array_muxed0 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed0 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed0 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed0 <= 10'd683;
		end
	endcase
// synthesis translate_off
	dummy_d_210 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_211;
// synthesis translate_on
always @(*) begin
	sync_f_array_muxed1 <= 10'd0;
	case (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c2)
		1'd0: begin
			sync_f_array_muxed1 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed1 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed1 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed1 <= 10'd683;
		end
	endcase
// synthesis translate_off
	dummy_d_211 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_212;
// synthesis translate_on
always @(*) begin
	sync_f_array_muxed2 <= 10'd0;
	case (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c2)
		1'd0: begin
			sync_f_array_muxed2 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed2 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed2 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed2 <= 10'd683;
		end
	endcase
// synthesis translate_off
	dummy_d_212 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_213;
// synthesis translate_on
always @(*) begin
	sync_f_array_muxed3 <= 10'd0;
	case (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c2)
		1'd0: begin
			sync_f_array_muxed3 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed3 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed3 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed3 <= 10'd683;
		end
	endcase
// synthesis translate_off
	dummy_d_213 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_214;
// synthesis translate_on
always @(*) begin
	sync_f_array_muxed4 <= 10'd0;
	case (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c2)
		1'd0: begin
			sync_f_array_muxed4 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed4 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed4 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed4 <= 10'd683;
		end
	endcase
// synthesis translate_off
	dummy_d_214 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_215;
// synthesis translate_on
always @(*) begin
	sync_f_array_muxed5 <= 10'd0;
	case (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c2)
		1'd0: begin
			sync_f_array_muxed5 <= 10'd852;
		end
		1'd1: begin
			sync_f_array_muxed5 <= 8'd171;
		end
		2'd2: begin
			sync_f_array_muxed5 <= 9'd340;
		end
		default: begin
			sync_f_array_muxed5 <= 10'd683;
		end
	endcase
// synthesis translate_off
	dummy_d_215 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_216;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed0 <= 13'd0;
	case (hdmi2usbsoc_ddrphy_phase_sel)
		1'd0: begin
			sync_rhs_array_muxed0 <= hdmi2usbsoc_ddrphy_record0_address;
		end
		default: begin
			sync_rhs_array_muxed0 <= hdmi2usbsoc_ddrphy_record1_address;
		end
	endcase
// synthesis translate_off
	dummy_d_216 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_217;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed1 <= 3'd0;
	case (hdmi2usbsoc_ddrphy_phase_sel)
		1'd0: begin
			sync_rhs_array_muxed1 <= hdmi2usbsoc_ddrphy_record0_bank;
		end
		default: begin
			sync_rhs_array_muxed1 <= hdmi2usbsoc_ddrphy_record1_bank;
		end
	endcase
// synthesis translate_off
	dummy_d_217 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_218;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed2 <= 1'd0;
	case (hdmi2usbsoc_ddrphy_phase_sel)
		1'd0: begin
			sync_rhs_array_muxed2 <= hdmi2usbsoc_ddrphy_record0_cke;
		end
		default: begin
			sync_rhs_array_muxed2 <= hdmi2usbsoc_ddrphy_record1_cke;
		end
	endcase
// synthesis translate_off
	dummy_d_218 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_219;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed3 <= 1'd0;
	case (hdmi2usbsoc_ddrphy_phase_sel)
		1'd0: begin
			sync_rhs_array_muxed3 <= hdmi2usbsoc_ddrphy_record0_ras_n;
		end
		default: begin
			sync_rhs_array_muxed3 <= hdmi2usbsoc_ddrphy_record1_ras_n;
		end
	endcase
// synthesis translate_off
	dummy_d_219 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_220;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed4 <= 1'd0;
	case (hdmi2usbsoc_ddrphy_phase_sel)
		1'd0: begin
			sync_rhs_array_muxed4 <= hdmi2usbsoc_ddrphy_record0_cas_n;
		end
		default: begin
			sync_rhs_array_muxed4 <= hdmi2usbsoc_ddrphy_record1_cas_n;
		end
	endcase
// synthesis translate_off
	dummy_d_220 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_221;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed5 <= 1'd0;
	case (hdmi2usbsoc_ddrphy_phase_sel)
		1'd0: begin
			sync_rhs_array_muxed5 <= hdmi2usbsoc_ddrphy_record0_we_n;
		end
		default: begin
			sync_rhs_array_muxed5 <= hdmi2usbsoc_ddrphy_record1_we_n;
		end
	endcase
// synthesis translate_off
	dummy_d_221 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_222;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed6 <= 1'd0;
	case (hdmi2usbsoc_ddrphy_phase_sel)
		1'd0: begin
			sync_rhs_array_muxed6 <= hdmi2usbsoc_ddrphy_record0_odt;
		end
		default: begin
			sync_rhs_array_muxed6 <= hdmi2usbsoc_ddrphy_record1_odt;
		end
	endcase
// synthesis translate_off
	dummy_d_222 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_223;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed7 <= 13'd0;
	case (hdmi2usbsoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed7 <= hdmi2usbsoc_sdram_nop_a;
		end
		1'd1: begin
			sync_rhs_array_muxed7 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			sync_rhs_array_muxed7 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			sync_rhs_array_muxed7 <= hdmi2usbsoc_sdram_cmd_payload_a;
		end
	endcase
// synthesis translate_off
	dummy_d_223 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_224;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed8 <= 3'd0;
	case (hdmi2usbsoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed8 <= hdmi2usbsoc_sdram_nop_ba;
		end
		1'd1: begin
			sync_rhs_array_muxed8 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			sync_rhs_array_muxed8 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			sync_rhs_array_muxed8 <= hdmi2usbsoc_sdram_cmd_payload_ba;
		end
	endcase
// synthesis translate_off
	dummy_d_224 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_225;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed9 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed9 <= hdmi2usbsoc_sdram_nop_cas;
		end
		1'd1: begin
			sync_rhs_array_muxed9 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			sync_rhs_array_muxed9 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			sync_rhs_array_muxed9 <= hdmi2usbsoc_sdram_cmd_payload_cas;
		end
	endcase
// synthesis translate_off
	dummy_d_225 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_226;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed10 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed10 <= hdmi2usbsoc_sdram_nop_ras;
		end
		1'd1: begin
			sync_rhs_array_muxed10 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			sync_rhs_array_muxed10 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			sync_rhs_array_muxed10 <= hdmi2usbsoc_sdram_cmd_payload_ras;
		end
	endcase
// synthesis translate_off
	dummy_d_226 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_227;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed11 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed11 <= hdmi2usbsoc_sdram_nop_we;
		end
		1'd1: begin
			sync_rhs_array_muxed11 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			sync_rhs_array_muxed11 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			sync_rhs_array_muxed11 <= hdmi2usbsoc_sdram_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_227 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_228;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed12 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed12 <= (hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			sync_rhs_array_muxed12 <= (hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			sync_rhs_array_muxed12 <= (hdmi2usbsoc_sdram_cmd_valid & hdmi2usbsoc_sdram_cmd_payload_is_read);
		end
	endcase
// synthesis translate_off
	dummy_d_228 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_229;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed13 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel0)
		1'd0: begin
			sync_rhs_array_muxed13 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed13 <= (hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			sync_rhs_array_muxed13 <= (hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			sync_rhs_array_muxed13 <= (hdmi2usbsoc_sdram_cmd_valid & hdmi2usbsoc_sdram_cmd_payload_is_write);
		end
	endcase
// synthesis translate_off
	dummy_d_229 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_230;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed14 <= 13'd0;
	case (hdmi2usbsoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed14 <= hdmi2usbsoc_sdram_nop_a;
		end
		1'd1: begin
			sync_rhs_array_muxed14 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			sync_rhs_array_muxed14 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			sync_rhs_array_muxed14 <= hdmi2usbsoc_sdram_cmd_payload_a;
		end
	endcase
// synthesis translate_off
	dummy_d_230 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_231;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed15 <= 3'd0;
	case (hdmi2usbsoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed15 <= hdmi2usbsoc_sdram_nop_ba;
		end
		1'd1: begin
			sync_rhs_array_muxed15 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			sync_rhs_array_muxed15 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			sync_rhs_array_muxed15 <= hdmi2usbsoc_sdram_cmd_payload_ba;
		end
	endcase
// synthesis translate_off
	dummy_d_231 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_232;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed16 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed16 <= hdmi2usbsoc_sdram_nop_cas;
		end
		1'd1: begin
			sync_rhs_array_muxed16 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			sync_rhs_array_muxed16 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			sync_rhs_array_muxed16 <= hdmi2usbsoc_sdram_cmd_payload_cas;
		end
	endcase
// synthesis translate_off
	dummy_d_232 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_233;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed17 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed17 <= hdmi2usbsoc_sdram_nop_ras;
		end
		1'd1: begin
			sync_rhs_array_muxed17 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			sync_rhs_array_muxed17 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			sync_rhs_array_muxed17 <= hdmi2usbsoc_sdram_cmd_payload_ras;
		end
	endcase
// synthesis translate_off
	dummy_d_233 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_234;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed18 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed18 <= hdmi2usbsoc_sdram_nop_we;
		end
		1'd1: begin
			sync_rhs_array_muxed18 <= hdmi2usbsoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			sync_rhs_array_muxed18 <= hdmi2usbsoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			sync_rhs_array_muxed18 <= hdmi2usbsoc_sdram_cmd_payload_we;
		end
	endcase
// synthesis translate_off
	dummy_d_234 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_235;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed19 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed19 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed19 <= (hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			sync_rhs_array_muxed19 <= (hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			sync_rhs_array_muxed19 <= (hdmi2usbsoc_sdram_cmd_valid & hdmi2usbsoc_sdram_cmd_payload_is_read);
		end
	endcase
// synthesis translate_off
	dummy_d_235 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_236;
// synthesis translate_on
always @(*) begin
	sync_rhs_array_muxed20 <= 1'd0;
	case (hdmi2usbsoc_sdram_sel1)
		1'd0: begin
			sync_rhs_array_muxed20 <= 1'd0;
		end
		1'd1: begin
			sync_rhs_array_muxed20 <= (hdmi2usbsoc_sdram_choose_cmd_cmd_valid & hdmi2usbsoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			sync_rhs_array_muxed20 <= (hdmi2usbsoc_sdram_choose_req_cmd_valid & hdmi2usbsoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			sync_rhs_array_muxed20 <= (hdmi2usbsoc_sdram_cmd_valid & hdmi2usbsoc_sdram_cmd_payload_is_write);
		end
	endcase
// synthesis translate_off
	dummy_d_236 <= dummy_s;
// synthesis translate_on
end
assign hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx = xilinxmultiregimpl0_regs1;
assign xilinxasyncresetsynchronizerimpl0 = ((~cpu_reset) | hdmi2usbsoc_crg_reset);
assign xilinxasyncresetsynchronizerimpl1 = ((~hdmi2usbsoc_crg_pll_lckd) | (hdmi2usbsoc_crg_por > 1'd0));
assign xilinxasyncresetsynchronizerimpl2 = (sys_rst | (~hdmi2usbsoc_crg_dcm_base50_locked));
assign hdmi2usbsoc_hdmi_in0_edid_scl_raw = xilinxmultiregimpl1_regs1;
assign hdmi2usbsoc_hdmi_in0_edid_sda_raw = xilinxmultiregimpl2_regs1;
assign hdmi2usbsoc_hdmi_in0_locked = xilinxmultiregimpl3_regs1;
assign xilinxasyncresetsynchronizerimpl4 = (~hdmi2usbsoc_hdmi_in0_locked_async);
assign xilinxasyncresetsynchronizerimpl5 = (~hdmi2usbsoc_hdmi_in0_locked_async);
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_o = xilinxmultiregimpl4_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_o = xilinxmultiregimpl5_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_o = xilinxmultiregimpl6_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_o = xilinxmultiregimpl7_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_o = xilinxmultiregimpl8_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_o = xilinxmultiregimpl9_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_o = xilinxmultiregimpl10_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_o = xilinxmultiregimpl11_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_status = xilinxmultiregimpl12_regs1;
assign xilinxmultiregimpl12 = {hdmi2usbsoc_hdmi_in0_s6datacapture0_too_early, hdmi2usbsoc_hdmi_in0_s6datacapture0_too_late};
assign hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_o = xilinxmultiregimpl13_regs1;
assign hdmi2usbsoc_hdmi_in0_charsync0_char_synced_status = xilinxmultiregimpl14_regs1;
assign hdmi2usbsoc_hdmi_in0_charsync0_ctl_pos_status = xilinxmultiregimpl15_regs1;
assign hdmi2usbsoc_hdmi_in0_wer0_toggle_o = xilinxmultiregimpl16_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_o = xilinxmultiregimpl17_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_o = xilinxmultiregimpl18_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_o = xilinxmultiregimpl19_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_o = xilinxmultiregimpl20_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_o = xilinxmultiregimpl21_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_o = xilinxmultiregimpl22_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_o = xilinxmultiregimpl23_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_o = xilinxmultiregimpl24_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_status = xilinxmultiregimpl25_regs1;
assign xilinxmultiregimpl25 = {hdmi2usbsoc_hdmi_in0_s6datacapture1_too_early, hdmi2usbsoc_hdmi_in0_s6datacapture1_too_late};
assign hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_o = xilinxmultiregimpl26_regs1;
assign hdmi2usbsoc_hdmi_in0_charsync1_char_synced_status = xilinxmultiregimpl27_regs1;
assign hdmi2usbsoc_hdmi_in0_charsync1_ctl_pos_status = xilinxmultiregimpl28_regs1;
assign hdmi2usbsoc_hdmi_in0_wer1_toggle_o = xilinxmultiregimpl29_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_o = xilinxmultiregimpl30_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_o = xilinxmultiregimpl31_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_o = xilinxmultiregimpl32_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_o = xilinxmultiregimpl33_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_o = xilinxmultiregimpl34_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_o = xilinxmultiregimpl35_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_o = xilinxmultiregimpl36_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_o = xilinxmultiregimpl37_regs1;
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_status = xilinxmultiregimpl38_regs1;
assign xilinxmultiregimpl38 = {hdmi2usbsoc_hdmi_in0_s6datacapture2_too_early, hdmi2usbsoc_hdmi_in0_s6datacapture2_too_late};
assign hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_o = xilinxmultiregimpl39_regs1;
assign hdmi2usbsoc_hdmi_in0_charsync2_char_synced_status = xilinxmultiregimpl40_regs1;
assign hdmi2usbsoc_hdmi_in0_charsync2_ctl_pos_status = xilinxmultiregimpl41_regs1;
assign hdmi2usbsoc_hdmi_in0_wer2_toggle_o = xilinxmultiregimpl42_regs1;
assign hdmi2usbsoc_hdmi_in0_chansync_status = xilinxmultiregimpl43_regs1;
assign hdmi2usbsoc_hdmi_in0_resdetection_hres_status = xilinxmultiregimpl44_regs1;
assign hdmi2usbsoc_hdmi_in0_resdetection_vres_status = xilinxmultiregimpl45_regs1;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_produce_rdomain = xilinxmultiregimpl46_regs1;
assign hdmi2usbsoc_hdmi_in0_frame_fifo_consume_wdomain = xilinxmultiregimpl47_regs1;
assign hdmi2usbsoc_hdmi_in0_frame_sys_overflow = xilinxmultiregimpl48_regs1;
assign hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_o = xilinxmultiregimpl49_regs1;
assign hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_o = xilinxmultiregimpl50_regs1;
assign hdmi2usbsoc_hdmi_in1_edid_scl_raw = xilinxmultiregimpl51_regs1;
assign hdmi2usbsoc_hdmi_in1_edid_sda_raw = xilinxmultiregimpl52_regs1;
assign hdmi2usbsoc_hdmi_in1_locked = xilinxmultiregimpl53_regs1;
assign xilinxasyncresetsynchronizerimpl6 = (~hdmi2usbsoc_hdmi_in1_locked_async);
assign xilinxasyncresetsynchronizerimpl7 = (~hdmi2usbsoc_hdmi_in1_locked_async);
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_o = xilinxmultiregimpl54_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_o = xilinxmultiregimpl55_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_o = xilinxmultiregimpl56_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_o = xilinxmultiregimpl57_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_o = xilinxmultiregimpl58_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_o = xilinxmultiregimpl59_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_o = xilinxmultiregimpl60_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_o = xilinxmultiregimpl61_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_status = xilinxmultiregimpl62_regs1;
assign xilinxmultiregimpl62 = {hdmi2usbsoc_hdmi_in1_s6datacapture0_too_early, hdmi2usbsoc_hdmi_in1_s6datacapture0_too_late};
assign hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_o = xilinxmultiregimpl63_regs1;
assign hdmi2usbsoc_hdmi_in1_charsync0_char_synced_status = xilinxmultiregimpl64_regs1;
assign hdmi2usbsoc_hdmi_in1_charsync0_ctl_pos_status = xilinxmultiregimpl65_regs1;
assign hdmi2usbsoc_hdmi_in1_wer0_toggle_o = xilinxmultiregimpl66_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_o = xilinxmultiregimpl67_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_o = xilinxmultiregimpl68_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_o = xilinxmultiregimpl69_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_o = xilinxmultiregimpl70_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_o = xilinxmultiregimpl71_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_o = xilinxmultiregimpl72_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_o = xilinxmultiregimpl73_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_o = xilinxmultiregimpl74_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_status = xilinxmultiregimpl75_regs1;
assign xilinxmultiregimpl75 = {hdmi2usbsoc_hdmi_in1_s6datacapture1_too_early, hdmi2usbsoc_hdmi_in1_s6datacapture1_too_late};
assign hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_o = xilinxmultiregimpl76_regs1;
assign hdmi2usbsoc_hdmi_in1_charsync1_char_synced_status = xilinxmultiregimpl77_regs1;
assign hdmi2usbsoc_hdmi_in1_charsync1_ctl_pos_status = xilinxmultiregimpl78_regs1;
assign hdmi2usbsoc_hdmi_in1_wer1_toggle_o = xilinxmultiregimpl79_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_o = xilinxmultiregimpl80_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_o = xilinxmultiregimpl81_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_o = xilinxmultiregimpl82_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_o = xilinxmultiregimpl83_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_o = xilinxmultiregimpl84_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_o = xilinxmultiregimpl85_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_o = xilinxmultiregimpl86_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_o = xilinxmultiregimpl87_regs1;
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_status = xilinxmultiregimpl88_regs1;
assign xilinxmultiregimpl88 = {hdmi2usbsoc_hdmi_in1_s6datacapture2_too_early, hdmi2usbsoc_hdmi_in1_s6datacapture2_too_late};
assign hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_o = xilinxmultiregimpl89_regs1;
assign hdmi2usbsoc_hdmi_in1_charsync2_char_synced_status = xilinxmultiregimpl90_regs1;
assign hdmi2usbsoc_hdmi_in1_charsync2_ctl_pos_status = xilinxmultiregimpl91_regs1;
assign hdmi2usbsoc_hdmi_in1_wer2_toggle_o = xilinxmultiregimpl92_regs1;
assign hdmi2usbsoc_hdmi_in1_chansync_status = xilinxmultiregimpl93_regs1;
assign hdmi2usbsoc_hdmi_in1_resdetection_hres_status = xilinxmultiregimpl94_regs1;
assign hdmi2usbsoc_hdmi_in1_resdetection_vres_status = xilinxmultiregimpl95_regs1;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_produce_rdomain = xilinxmultiregimpl96_regs1;
assign hdmi2usbsoc_hdmi_in1_frame_fifo_consume_wdomain = xilinxmultiregimpl97_regs1;
assign hdmi2usbsoc_hdmi_in1_frame_sys_overflow = xilinxmultiregimpl98_regs1;
assign hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_o = xilinxmultiregimpl99_regs1;
assign hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_o = xilinxmultiregimpl100_regs1;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_produce_rdomain = xilinxmultiregimpl101_regs1;
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_consume_wdomain = xilinxmultiregimpl102_regs1;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_produce_rdomain = xilinxmultiregimpl103_regs1;
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_consume_wdomain = xilinxmultiregimpl104_regs1;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_produce_rdomain = xilinxmultiregimpl105_regs1;
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_consume_wdomain = xilinxmultiregimpl106_regs1;
assign hdmi2usbsoc_hdmi_out0_core_underflow_enable = xilinxmultiregimpl107_regs1;
assign hdmi2usbsoc_hdmi_out0_core_toggle_o = xilinxmultiregimpl108_regs1;
assign hdmi2usbsoc_hdmi_out0_driver_clocking_mult_locked = xilinxmultiregimpl109_regs1;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_produce_rdomain = xilinxmultiregimpl110_regs1;
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_consume_wdomain = xilinxmultiregimpl111_regs1;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_produce_rdomain = xilinxmultiregimpl112_regs1;
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_consume_wdomain = xilinxmultiregimpl113_regs1;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_produce_rdomain = xilinxmultiregimpl114_regs1;
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_consume_wdomain = xilinxmultiregimpl115_regs1;
assign hdmi2usbsoc_hdmi_out1_core_underflow_enable = xilinxmultiregimpl116_regs1;
assign hdmi2usbsoc_hdmi_out1_core_toggle_o = xilinxmultiregimpl117_regs1;
assign encoder_cdc_produce_rdomain = xilinxmultiregimpl118_regs1;
assign encoder_cdc_consume_wdomain = xilinxmultiregimpl119_regs1;
assign encoder_streamer_fifo_produce_rdomain = xilinxmultiregimpl120_regs1;
assign encoder_streamer_fifo_consume_wdomain = xilinxmultiregimpl121_regs1;

always @(posedge encoder_clk) begin
	encoder_cdc_graycounter1_q_binary <= encoder_cdc_graycounter1_q_next_binary;
	encoder_cdc_graycounter1_q <= encoder_cdc_graycounter1_q_next;
	if (encoderbuffer_write_swap) begin
		encoderbuffer_write_sel <= (~encoderbuffer_write_sel);
	end
	if (encoderbuffer_read_swap) begin
		encoderbuffer_read_sel <= (~encoderbuffer_read_sel);
	end
	if (encoderbuffer_v_write_clr) begin
		encoderbuffer_v_write <= 1'd0;
	end else begin
		if (encoderbuffer_v_write_inc) begin
			encoderbuffer_v_write <= (encoderbuffer_v_write + 1'd1);
		end
	end
	if (encoderbuffer_h_read_clr) begin
		encoderbuffer_h_read <= 1'd0;
	end else begin
		if (encoderbuffer_h_read_inc) begin
			encoderbuffer_h_read <= (encoderbuffer_h_read + 1'd1);
		end
	end
	if (encoderbuffer_v_read_clr) begin
		encoderbuffer_v_read <= 1'd0;
	end else begin
		if (encoderbuffer_v_read_inc) begin
			encoderbuffer_v_read <= (encoderbuffer_v_read + 1'd1);
		end
	end
	fsm0_state <= fsm0_next_state;
	fsm1_state <= fsm1_next_state;
	if (encoder_fdct_fifo_rd) begin
		encoder_fdct_data_d1 <= {encoder_source_source_payload_cr, encoder_source_source_payload_cb, encoder_source_source_payload_y};
	end
	encoder_fdct_data_d2 <= encoder_fdct_data_d1;
	encoder_fdct_data_d3 <= encoder_fdct_data_d2;
	encoder_fdct_data_d4 <= encoder_fdct_data_d3;
	encoder_fdct_data_d5 <= encoder_fdct_data_d4;
	if ((encoder_sink_sink_valid1 & encoder_sink_sink_ready1)) begin
		encoder_parity_in <= (~encoder_parity_in);
	end
	if ((encoder_source_source_valid1 & encoder_source_source_ready1)) begin
		encoder_parity_out <= (~encoder_parity_out);
	end
	if (((encoder_y_fifo_syncfifo_we & encoder_y_fifo_syncfifo_writable) & (~encoder_y_fifo_replace))) begin
		encoder_y_fifo_produce <= (encoder_y_fifo_produce + 1'd1);
	end
	if (encoder_y_fifo_do_read) begin
		encoder_y_fifo_consume <= (encoder_y_fifo_consume + 1'd1);
	end
	if (((encoder_y_fifo_syncfifo_we & encoder_y_fifo_syncfifo_writable) & (~encoder_y_fifo_replace))) begin
		if ((~encoder_y_fifo_do_read)) begin
			encoder_y_fifo_level <= (encoder_y_fifo_level + 1'd1);
		end
	end else begin
		if (encoder_y_fifo_do_read) begin
			encoder_y_fifo_level <= (encoder_y_fifo_level - 1'd1);
		end
	end
	if (((encoder_cb_fifo_syncfifo_we & encoder_cb_fifo_syncfifo_writable) & (~encoder_cb_fifo_replace))) begin
		encoder_cb_fifo_produce <= (encoder_cb_fifo_produce + 1'd1);
	end
	if (encoder_cb_fifo_do_read) begin
		encoder_cb_fifo_consume <= (encoder_cb_fifo_consume + 1'd1);
	end
	if (((encoder_cb_fifo_syncfifo_we & encoder_cb_fifo_syncfifo_writable) & (~encoder_cb_fifo_replace))) begin
		if ((~encoder_cb_fifo_do_read)) begin
			encoder_cb_fifo_level <= (encoder_cb_fifo_level + 1'd1);
		end
	end else begin
		if (encoder_cb_fifo_do_read) begin
			encoder_cb_fifo_level <= (encoder_cb_fifo_level - 1'd1);
		end
	end
	if (((encoder_cr_fifo_syncfifo_we & encoder_cr_fifo_syncfifo_writable) & (~encoder_cr_fifo_replace))) begin
		encoder_cr_fifo_produce <= (encoder_cr_fifo_produce + 1'd1);
	end
	if (encoder_cr_fifo_do_read) begin
		encoder_cr_fifo_consume <= (encoder_cr_fifo_consume + 1'd1);
	end
	if (((encoder_cr_fifo_syncfifo_we & encoder_cr_fifo_syncfifo_writable) & (~encoder_cr_fifo_replace))) begin
		if ((~encoder_cr_fifo_do_read)) begin
			encoder_cr_fifo_level <= (encoder_cr_fifo_level + 1'd1);
		end
	end else begin
		if (encoder_cr_fifo_do_read) begin
			encoder_cr_fifo_level <= (encoder_cr_fifo_level - 1'd1);
		end
	end
	if (encoder_reset) begin
		encoder_y_fifo_level <= 3'd0;
		encoder_y_fifo_produce <= 2'd0;
		encoder_y_fifo_consume <= 2'd0;
		encoder_cb_fifo_level <= 3'd0;
		encoder_cb_fifo_produce <= 2'd0;
		encoder_cb_fifo_consume <= 2'd0;
		encoder_cr_fifo_level <= 3'd0;
		encoder_cr_fifo_produce <= 2'd0;
		encoder_cr_fifo_consume <= 2'd0;
		encoder_parity_in <= 1'd0;
		encoder_parity_out <= 1'd0;
	end
	if (encoder_output_fifo_syncfifo_re) begin
		encoder_output_fifo_readable <= 1'd1;
	end else begin
		if (encoder_output_fifo_re) begin
			encoder_output_fifo_readable <= 1'd0;
		end
	end
	if (((encoder_output_fifo_syncfifo_we & encoder_output_fifo_syncfifo_writable) & (~encoder_output_fifo_replace))) begin
		encoder_output_fifo_produce <= (encoder_output_fifo_produce + 1'd1);
	end
	if (encoder_output_fifo_do_read) begin
		encoder_output_fifo_consume <= (encoder_output_fifo_consume + 1'd1);
	end
	if (((encoder_output_fifo_syncfifo_we & encoder_output_fifo_syncfifo_writable) & (~encoder_output_fifo_replace))) begin
		if ((~encoder_output_fifo_do_read)) begin
			encoder_output_fifo_level0 <= (encoder_output_fifo_level0 + 1'd1);
		end
	end else begin
		if (encoder_output_fifo_do_read) begin
			encoder_output_fifo_level0 <= (encoder_output_fifo_level0 - 1'd1);
		end
	end
	encoder_streamer_fifo_graycounter0_q_binary <= encoder_streamer_fifo_graycounter0_q_next_binary;
	encoder_streamer_fifo_graycounter0_q <= encoder_streamer_fifo_graycounter0_q_next;
	if (encoder_rst) begin
		encoder_cdc_graycounter1_q <= 3'd0;
		encoder_cdc_graycounter1_q_binary <= 3'd0;
		encoderbuffer_write_sel <= 1'd0;
		encoderbuffer_read_sel <= 1'd1;
		encoderbuffer_v_write <= 3'd0;
		encoderbuffer_h_read <= 3'd0;
		encoderbuffer_v_read <= 3'd0;
		encoder_y_fifo_level <= 3'd0;
		encoder_y_fifo_produce <= 2'd0;
		encoder_y_fifo_consume <= 2'd0;
		encoder_cb_fifo_level <= 3'd0;
		encoder_cb_fifo_produce <= 2'd0;
		encoder_cb_fifo_consume <= 2'd0;
		encoder_cr_fifo_level <= 3'd0;
		encoder_cr_fifo_produce <= 2'd0;
		encoder_cr_fifo_consume <= 2'd0;
		encoder_parity_in <= 1'd0;
		encoder_parity_out <= 1'd0;
		encoder_fdct_data_d1 <= 24'd0;
		encoder_fdct_data_d2 <= 24'd0;
		encoder_fdct_data_d3 <= 24'd0;
		encoder_fdct_data_d4 <= 24'd0;
		encoder_fdct_data_d5 <= 24'd0;
		encoder_output_fifo_readable <= 1'd0;
		encoder_output_fifo_level0 <= 11'd0;
		encoder_output_fifo_produce <= 10'd0;
		encoder_output_fifo_consume <= 10'd0;
		encoder_streamer_fifo_graycounter0_q <= 3'd0;
		encoder_streamer_fifo_graycounter0_q_binary <= 3'd0;
		fsm0_state <= 1'd0;
		fsm1_state <= 1'd0;
	end
	xilinxmultiregimpl118_regs0 <= encoder_cdc_graycounter0_q;
	xilinxmultiregimpl118_regs1 <= xilinxmultiregimpl118_regs0;
	xilinxmultiregimpl121_regs0 <= encoder_streamer_fifo_graycounter1_q;
	xilinxmultiregimpl121_regs1 <= xilinxmultiregimpl121_regs0;
end

always @(posedge hdmi_in0_pix_clk) begin
	hdmi2usbsoc_hdmi_in0_s6datacapture0_d <= hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr;
	hdmi2usbsoc_hdmi_in0_charsync0_raw_data1 <= hdmi2usbsoc_hdmi_in0_charsync0_raw_data;
	hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd0;
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[9:0] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[9:0] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[9:0] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[9:0] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 1'd0;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[10:1] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[10:1] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[10:1] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[10:1] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 1'd1;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[11:2] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[11:2] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[11:2] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[11:2] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 2'd2;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[12:3] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[12:3] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[12:3] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[12:3] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 2'd3;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[13:4] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[13:4] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[13:4] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[13:4] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 3'd4;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[14:5] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[14:5] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[14:5] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[14:5] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 3'd5;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[15:6] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[15:6] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[15:6] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[15:6] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 3'd6;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[16:7] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[16:7] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[16:7] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[16:7] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 3'd7;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[17:8] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[17:8] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[17:8] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[17:8] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 4'd8;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync0_raw[18:9] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[18:9] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[18:9] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync0_raw[18:9] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 4'd9;
	end
	if ((hdmi2usbsoc_hdmi_in0_charsync0_found_control & (hdmi2usbsoc_hdmi_in0_charsync0_control_position == hdmi2usbsoc_hdmi_in0_charsync0_previous_control_position))) begin
		if ((hdmi2usbsoc_hdmi_in0_charsync0_control_counter == 3'd7)) begin
			hdmi2usbsoc_hdmi_in0_charsync0_control_counter <= 1'd0;
			hdmi2usbsoc_hdmi_in0_charsync0_synced <= 1'd1;
			hdmi2usbsoc_hdmi_in0_charsync0_word_sel <= hdmi2usbsoc_hdmi_in0_charsync0_control_position;
		end else begin
			hdmi2usbsoc_hdmi_in0_charsync0_control_counter <= (hdmi2usbsoc_hdmi_in0_charsync0_control_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_in0_charsync0_control_counter <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in0_charsync0_previous_control_position <= hdmi2usbsoc_hdmi_in0_charsync0_control_position;
	hdmi2usbsoc_hdmi_in0_charsync0_data <= (hdmi2usbsoc_hdmi_in0_charsync0_raw >>> hdmi2usbsoc_hdmi_in0_charsync0_word_sel);
	hdmi2usbsoc_hdmi_in0_wer0_data_r <= hdmi2usbsoc_hdmi_in0_wer0_data[8:0];
	hdmi2usbsoc_hdmi_in0_wer0_transition_count <= (((((((hdmi2usbsoc_hdmi_in0_wer0_transitions[0] + hdmi2usbsoc_hdmi_in0_wer0_transitions[1]) + hdmi2usbsoc_hdmi_in0_wer0_transitions[2]) + hdmi2usbsoc_hdmi_in0_wer0_transitions[3]) + hdmi2usbsoc_hdmi_in0_wer0_transitions[4]) + hdmi2usbsoc_hdmi_in0_wer0_transitions[5]) + hdmi2usbsoc_hdmi_in0_wer0_transitions[6]) + hdmi2usbsoc_hdmi_in0_wer0_transitions[7]);
	hdmi2usbsoc_hdmi_in0_wer0_is_control <= ((((hdmi2usbsoc_hdmi_in0_wer0_data_r == 10'd852) | (hdmi2usbsoc_hdmi_in0_wer0_data_r == 8'd171)) | (hdmi2usbsoc_hdmi_in0_wer0_data_r == 9'd340)) | (hdmi2usbsoc_hdmi_in0_wer0_data_r == 10'd683));
	hdmi2usbsoc_hdmi_in0_wer0_is_error <= ((hdmi2usbsoc_hdmi_in0_wer0_transition_count > 3'd4) & (~hdmi2usbsoc_hdmi_in0_wer0_is_control));
	{hdmi2usbsoc_hdmi_in0_wer0_period_done, hdmi2usbsoc_hdmi_in0_wer0_period_counter} <= (hdmi2usbsoc_hdmi_in0_wer0_period_counter + 1'd1);
	hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r_updated <= hdmi2usbsoc_hdmi_in0_wer0_period_done;
	if (hdmi2usbsoc_hdmi_in0_wer0_period_done) begin
		hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r <= hdmi2usbsoc_hdmi_in0_wer0_wer_counter;
		hdmi2usbsoc_hdmi_in0_wer0_wer_counter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_wer0_is_error) begin
			hdmi2usbsoc_hdmi_in0_wer0_wer_counter <= (hdmi2usbsoc_hdmi_in0_wer0_wer_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in0_wer0_i) begin
		hdmi2usbsoc_hdmi_in0_wer0_toggle_i <= (~hdmi2usbsoc_hdmi_in0_wer0_toggle_i);
	end
	hdmi2usbsoc_hdmi_in0_decoding0_output_de <= 1'd1;
	if ((hdmi2usbsoc_hdmi_in0_decoding0_input == 10'd852)) begin
		hdmi2usbsoc_hdmi_in0_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_c <= 1'd0;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding0_input == 8'd171)) begin
		hdmi2usbsoc_hdmi_in0_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_c <= 1'd1;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding0_input == 9'd340)) begin
		hdmi2usbsoc_hdmi_in0_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_c <= 2'd2;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding0_input == 10'd683)) begin
		hdmi2usbsoc_hdmi_in0_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_c <= 2'd3;
	end
	hdmi2usbsoc_hdmi_in0_decoding0_output_raw <= hdmi2usbsoc_hdmi_in0_decoding0_input;
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[0] <= (hdmi2usbsoc_hdmi_in0_decoding0_input[0] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[9]);
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[1] <= ((hdmi2usbsoc_hdmi_in0_decoding0_input[1] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[0]) ^ (~hdmi2usbsoc_hdmi_in0_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[2] <= ((hdmi2usbsoc_hdmi_in0_decoding0_input[2] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[1]) ^ (~hdmi2usbsoc_hdmi_in0_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[3] <= ((hdmi2usbsoc_hdmi_in0_decoding0_input[3] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[2]) ^ (~hdmi2usbsoc_hdmi_in0_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[4] <= ((hdmi2usbsoc_hdmi_in0_decoding0_input[4] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[3]) ^ (~hdmi2usbsoc_hdmi_in0_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[5] <= ((hdmi2usbsoc_hdmi_in0_decoding0_input[5] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[4]) ^ (~hdmi2usbsoc_hdmi_in0_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[6] <= ((hdmi2usbsoc_hdmi_in0_decoding0_input[6] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[5]) ^ (~hdmi2usbsoc_hdmi_in0_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding0_output_d[7] <= ((hdmi2usbsoc_hdmi_in0_decoding0_input[7] ^ hdmi2usbsoc_hdmi_in0_decoding0_input[6]) ^ (~hdmi2usbsoc_hdmi_in0_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding0_valid_o <= hdmi2usbsoc_hdmi_in0_decoding0_valid_i;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_d <= hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr;
	hdmi2usbsoc_hdmi_in0_charsync1_raw_data1 <= hdmi2usbsoc_hdmi_in0_charsync1_raw_data;
	hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd0;
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[9:0] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[9:0] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[9:0] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[9:0] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 1'd0;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[10:1] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[10:1] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[10:1] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[10:1] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 1'd1;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[11:2] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[11:2] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[11:2] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[11:2] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 2'd2;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[12:3] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[12:3] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[12:3] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[12:3] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 2'd3;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[13:4] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[13:4] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[13:4] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[13:4] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 3'd4;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[14:5] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[14:5] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[14:5] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[14:5] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 3'd5;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[15:6] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[15:6] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[15:6] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[15:6] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 3'd6;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[16:7] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[16:7] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[16:7] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[16:7] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 3'd7;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[17:8] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[17:8] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[17:8] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[17:8] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 4'd8;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync1_raw[18:9] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[18:9] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[18:9] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync1_raw[18:9] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 4'd9;
	end
	if ((hdmi2usbsoc_hdmi_in0_charsync1_found_control & (hdmi2usbsoc_hdmi_in0_charsync1_control_position == hdmi2usbsoc_hdmi_in0_charsync1_previous_control_position))) begin
		if ((hdmi2usbsoc_hdmi_in0_charsync1_control_counter == 3'd7)) begin
			hdmi2usbsoc_hdmi_in0_charsync1_control_counter <= 1'd0;
			hdmi2usbsoc_hdmi_in0_charsync1_synced <= 1'd1;
			hdmi2usbsoc_hdmi_in0_charsync1_word_sel <= hdmi2usbsoc_hdmi_in0_charsync1_control_position;
		end else begin
			hdmi2usbsoc_hdmi_in0_charsync1_control_counter <= (hdmi2usbsoc_hdmi_in0_charsync1_control_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_in0_charsync1_control_counter <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in0_charsync1_previous_control_position <= hdmi2usbsoc_hdmi_in0_charsync1_control_position;
	hdmi2usbsoc_hdmi_in0_charsync1_data <= (hdmi2usbsoc_hdmi_in0_charsync1_raw >>> hdmi2usbsoc_hdmi_in0_charsync1_word_sel);
	hdmi2usbsoc_hdmi_in0_wer1_data_r <= hdmi2usbsoc_hdmi_in0_wer1_data[8:0];
	hdmi2usbsoc_hdmi_in0_wer1_transition_count <= (((((((hdmi2usbsoc_hdmi_in0_wer1_transitions[0] + hdmi2usbsoc_hdmi_in0_wer1_transitions[1]) + hdmi2usbsoc_hdmi_in0_wer1_transitions[2]) + hdmi2usbsoc_hdmi_in0_wer1_transitions[3]) + hdmi2usbsoc_hdmi_in0_wer1_transitions[4]) + hdmi2usbsoc_hdmi_in0_wer1_transitions[5]) + hdmi2usbsoc_hdmi_in0_wer1_transitions[6]) + hdmi2usbsoc_hdmi_in0_wer1_transitions[7]);
	hdmi2usbsoc_hdmi_in0_wer1_is_control <= ((((hdmi2usbsoc_hdmi_in0_wer1_data_r == 10'd852) | (hdmi2usbsoc_hdmi_in0_wer1_data_r == 8'd171)) | (hdmi2usbsoc_hdmi_in0_wer1_data_r == 9'd340)) | (hdmi2usbsoc_hdmi_in0_wer1_data_r == 10'd683));
	hdmi2usbsoc_hdmi_in0_wer1_is_error <= ((hdmi2usbsoc_hdmi_in0_wer1_transition_count > 3'd4) & (~hdmi2usbsoc_hdmi_in0_wer1_is_control));
	{hdmi2usbsoc_hdmi_in0_wer1_period_done, hdmi2usbsoc_hdmi_in0_wer1_period_counter} <= (hdmi2usbsoc_hdmi_in0_wer1_period_counter + 1'd1);
	hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r_updated <= hdmi2usbsoc_hdmi_in0_wer1_period_done;
	if (hdmi2usbsoc_hdmi_in0_wer1_period_done) begin
		hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r <= hdmi2usbsoc_hdmi_in0_wer1_wer_counter;
		hdmi2usbsoc_hdmi_in0_wer1_wer_counter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_wer1_is_error) begin
			hdmi2usbsoc_hdmi_in0_wer1_wer_counter <= (hdmi2usbsoc_hdmi_in0_wer1_wer_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in0_wer1_i) begin
		hdmi2usbsoc_hdmi_in0_wer1_toggle_i <= (~hdmi2usbsoc_hdmi_in0_wer1_toggle_i);
	end
	hdmi2usbsoc_hdmi_in0_decoding1_output_de <= 1'd1;
	if ((hdmi2usbsoc_hdmi_in0_decoding1_input == 10'd852)) begin
		hdmi2usbsoc_hdmi_in0_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_c <= 1'd0;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding1_input == 8'd171)) begin
		hdmi2usbsoc_hdmi_in0_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_c <= 1'd1;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding1_input == 9'd340)) begin
		hdmi2usbsoc_hdmi_in0_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_c <= 2'd2;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding1_input == 10'd683)) begin
		hdmi2usbsoc_hdmi_in0_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_c <= 2'd3;
	end
	hdmi2usbsoc_hdmi_in0_decoding1_output_raw <= hdmi2usbsoc_hdmi_in0_decoding1_input;
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[0] <= (hdmi2usbsoc_hdmi_in0_decoding1_input[0] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[9]);
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[1] <= ((hdmi2usbsoc_hdmi_in0_decoding1_input[1] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[0]) ^ (~hdmi2usbsoc_hdmi_in0_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[2] <= ((hdmi2usbsoc_hdmi_in0_decoding1_input[2] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[1]) ^ (~hdmi2usbsoc_hdmi_in0_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[3] <= ((hdmi2usbsoc_hdmi_in0_decoding1_input[3] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[2]) ^ (~hdmi2usbsoc_hdmi_in0_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[4] <= ((hdmi2usbsoc_hdmi_in0_decoding1_input[4] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[3]) ^ (~hdmi2usbsoc_hdmi_in0_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[5] <= ((hdmi2usbsoc_hdmi_in0_decoding1_input[5] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[4]) ^ (~hdmi2usbsoc_hdmi_in0_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[6] <= ((hdmi2usbsoc_hdmi_in0_decoding1_input[6] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[5]) ^ (~hdmi2usbsoc_hdmi_in0_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding1_output_d[7] <= ((hdmi2usbsoc_hdmi_in0_decoding1_input[7] ^ hdmi2usbsoc_hdmi_in0_decoding1_input[6]) ^ (~hdmi2usbsoc_hdmi_in0_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding1_valid_o <= hdmi2usbsoc_hdmi_in0_decoding1_valid_i;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_d <= hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr;
	hdmi2usbsoc_hdmi_in0_charsync2_raw_data1 <= hdmi2usbsoc_hdmi_in0_charsync2_raw_data;
	hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd0;
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[9:0] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[9:0] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[9:0] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[9:0] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 1'd0;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[10:1] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[10:1] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[10:1] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[10:1] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 1'd1;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[11:2] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[11:2] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[11:2] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[11:2] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 2'd2;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[12:3] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[12:3] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[12:3] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[12:3] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 2'd3;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[13:4] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[13:4] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[13:4] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[13:4] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 3'd4;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[14:5] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[14:5] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[14:5] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[14:5] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 3'd5;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[15:6] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[15:6] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[15:6] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[15:6] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 3'd6;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[16:7] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[16:7] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[16:7] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[16:7] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 3'd7;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[17:8] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[17:8] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[17:8] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[17:8] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 4'd8;
	end
	if (((((hdmi2usbsoc_hdmi_in0_charsync2_raw[18:9] == 10'd852) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[18:9] == 8'd171)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[18:9] == 9'd340)) | (hdmi2usbsoc_hdmi_in0_charsync2_raw[18:9] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 4'd9;
	end
	if ((hdmi2usbsoc_hdmi_in0_charsync2_found_control & (hdmi2usbsoc_hdmi_in0_charsync2_control_position == hdmi2usbsoc_hdmi_in0_charsync2_previous_control_position))) begin
		if ((hdmi2usbsoc_hdmi_in0_charsync2_control_counter == 3'd7)) begin
			hdmi2usbsoc_hdmi_in0_charsync2_control_counter <= 1'd0;
			hdmi2usbsoc_hdmi_in0_charsync2_synced <= 1'd1;
			hdmi2usbsoc_hdmi_in0_charsync2_word_sel <= hdmi2usbsoc_hdmi_in0_charsync2_control_position;
		end else begin
			hdmi2usbsoc_hdmi_in0_charsync2_control_counter <= (hdmi2usbsoc_hdmi_in0_charsync2_control_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_in0_charsync2_control_counter <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in0_charsync2_previous_control_position <= hdmi2usbsoc_hdmi_in0_charsync2_control_position;
	hdmi2usbsoc_hdmi_in0_charsync2_data <= (hdmi2usbsoc_hdmi_in0_charsync2_raw >>> hdmi2usbsoc_hdmi_in0_charsync2_word_sel);
	hdmi2usbsoc_hdmi_in0_wer2_data_r <= hdmi2usbsoc_hdmi_in0_wer2_data[8:0];
	hdmi2usbsoc_hdmi_in0_wer2_transition_count <= (((((((hdmi2usbsoc_hdmi_in0_wer2_transitions[0] + hdmi2usbsoc_hdmi_in0_wer2_transitions[1]) + hdmi2usbsoc_hdmi_in0_wer2_transitions[2]) + hdmi2usbsoc_hdmi_in0_wer2_transitions[3]) + hdmi2usbsoc_hdmi_in0_wer2_transitions[4]) + hdmi2usbsoc_hdmi_in0_wer2_transitions[5]) + hdmi2usbsoc_hdmi_in0_wer2_transitions[6]) + hdmi2usbsoc_hdmi_in0_wer2_transitions[7]);
	hdmi2usbsoc_hdmi_in0_wer2_is_control <= ((((hdmi2usbsoc_hdmi_in0_wer2_data_r == 10'd852) | (hdmi2usbsoc_hdmi_in0_wer2_data_r == 8'd171)) | (hdmi2usbsoc_hdmi_in0_wer2_data_r == 9'd340)) | (hdmi2usbsoc_hdmi_in0_wer2_data_r == 10'd683));
	hdmi2usbsoc_hdmi_in0_wer2_is_error <= ((hdmi2usbsoc_hdmi_in0_wer2_transition_count > 3'd4) & (~hdmi2usbsoc_hdmi_in0_wer2_is_control));
	{hdmi2usbsoc_hdmi_in0_wer2_period_done, hdmi2usbsoc_hdmi_in0_wer2_period_counter} <= (hdmi2usbsoc_hdmi_in0_wer2_period_counter + 1'd1);
	hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r_updated <= hdmi2usbsoc_hdmi_in0_wer2_period_done;
	if (hdmi2usbsoc_hdmi_in0_wer2_period_done) begin
		hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r <= hdmi2usbsoc_hdmi_in0_wer2_wer_counter;
		hdmi2usbsoc_hdmi_in0_wer2_wer_counter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_wer2_is_error) begin
			hdmi2usbsoc_hdmi_in0_wer2_wer_counter <= (hdmi2usbsoc_hdmi_in0_wer2_wer_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in0_wer2_i) begin
		hdmi2usbsoc_hdmi_in0_wer2_toggle_i <= (~hdmi2usbsoc_hdmi_in0_wer2_toggle_i);
	end
	hdmi2usbsoc_hdmi_in0_decoding2_output_de <= 1'd1;
	if ((hdmi2usbsoc_hdmi_in0_decoding2_input == 10'd852)) begin
		hdmi2usbsoc_hdmi_in0_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_c <= 1'd0;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding2_input == 8'd171)) begin
		hdmi2usbsoc_hdmi_in0_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_c <= 1'd1;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding2_input == 9'd340)) begin
		hdmi2usbsoc_hdmi_in0_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_c <= 2'd2;
	end
	if ((hdmi2usbsoc_hdmi_in0_decoding2_input == 10'd683)) begin
		hdmi2usbsoc_hdmi_in0_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_c <= 2'd3;
	end
	hdmi2usbsoc_hdmi_in0_decoding2_output_raw <= hdmi2usbsoc_hdmi_in0_decoding2_input;
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[0] <= (hdmi2usbsoc_hdmi_in0_decoding2_input[0] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[9]);
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[1] <= ((hdmi2usbsoc_hdmi_in0_decoding2_input[1] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[0]) ^ (~hdmi2usbsoc_hdmi_in0_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[2] <= ((hdmi2usbsoc_hdmi_in0_decoding2_input[2] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[1]) ^ (~hdmi2usbsoc_hdmi_in0_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[3] <= ((hdmi2usbsoc_hdmi_in0_decoding2_input[3] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[2]) ^ (~hdmi2usbsoc_hdmi_in0_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[4] <= ((hdmi2usbsoc_hdmi_in0_decoding2_input[4] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[3]) ^ (~hdmi2usbsoc_hdmi_in0_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[5] <= ((hdmi2usbsoc_hdmi_in0_decoding2_input[5] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[4]) ^ (~hdmi2usbsoc_hdmi_in0_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[6] <= ((hdmi2usbsoc_hdmi_in0_decoding2_input[6] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[5]) ^ (~hdmi2usbsoc_hdmi_in0_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding2_output_d[7] <= ((hdmi2usbsoc_hdmi_in0_decoding2_input[7] ^ hdmi2usbsoc_hdmi_in0_decoding2_input[6]) ^ (~hdmi2usbsoc_hdmi_in0_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in0_decoding2_valid_o <= hdmi2usbsoc_hdmi_in0_decoding2_valid_i;
	if ((~hdmi2usbsoc_hdmi_in0_chansync_valid_i)) begin
		hdmi2usbsoc_hdmi_in0_chansync_chan_synced <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_chansync_some_control) begin
			if (hdmi2usbsoc_hdmi_in0_chansync_all_control) begin
				hdmi2usbsoc_hdmi_in0_chansync_chan_synced <= 1'd1;
			end else begin
				hdmi2usbsoc_hdmi_in0_chansync_chan_synced <= 1'd0;
			end
		end
	end
	hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_produce <= (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_produce + 1'd1);
	if (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_re) begin
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_consume <= (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_consume + 1'd1);
	end
	hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_produce <= (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_produce + 1'd1);
	if (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_re) begin
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_consume <= (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_consume + 1'd1);
	end
	hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_produce <= (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_produce + 1'd1);
	if (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_re) begin
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_consume <= (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_consume + 1'd1);
	end
	hdmi2usbsoc_hdmi_in0_syncpol_valid_o <= hdmi2usbsoc_hdmi_in0_syncpol_valid_i;
	hdmi2usbsoc_hdmi_in0_syncpol_r <= hdmi2usbsoc_hdmi_in0_syncpol_data_in2_d;
	hdmi2usbsoc_hdmi_in0_syncpol_g <= hdmi2usbsoc_hdmi_in0_syncpol_data_in1_d;
	hdmi2usbsoc_hdmi_in0_syncpol_b <= hdmi2usbsoc_hdmi_in0_syncpol_data_in0_d;
	hdmi2usbsoc_hdmi_in0_syncpol_de_r <= hdmi2usbsoc_hdmi_in0_syncpol_data_in0_de;
	if ((hdmi2usbsoc_hdmi_in0_syncpol_de_r & (~hdmi2usbsoc_hdmi_in0_syncpol_data_in0_de))) begin
		hdmi2usbsoc_hdmi_in0_syncpol_c_polarity <= hdmi2usbsoc_hdmi_in0_syncpol_data_in0_c;
		hdmi2usbsoc_hdmi_in0_syncpol_c_out <= 1'd0;
	end else begin
		hdmi2usbsoc_hdmi_in0_syncpol_c_out <= (hdmi2usbsoc_hdmi_in0_syncpol_data_in0_c ^ hdmi2usbsoc_hdmi_in0_syncpol_c_polarity);
	end
	hdmi2usbsoc_hdmi_in0_resdetection_de_r <= hdmi2usbsoc_hdmi_in0_resdetection_de;
	if ((hdmi2usbsoc_hdmi_in0_resdetection_valid_i & hdmi2usbsoc_hdmi_in0_resdetection_de)) begin
		hdmi2usbsoc_hdmi_in0_resdetection_hcounter <= (hdmi2usbsoc_hdmi_in0_resdetection_hcounter + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in0_resdetection_hcounter <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_in0_resdetection_valid_i) begin
		if (hdmi2usbsoc_hdmi_in0_resdetection_pn_de) begin
			hdmi2usbsoc_hdmi_in0_resdetection_hcounter_st <= hdmi2usbsoc_hdmi_in0_resdetection_hcounter;
		end
	end else begin
		hdmi2usbsoc_hdmi_in0_resdetection_hcounter_st <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in0_resdetection_vsync_r <= hdmi2usbsoc_hdmi_in0_resdetection_vsync;
	if ((hdmi2usbsoc_hdmi_in0_resdetection_valid_i & hdmi2usbsoc_hdmi_in0_resdetection_p_vsync)) begin
		hdmi2usbsoc_hdmi_in0_resdetection_vcounter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_resdetection_pn_de) begin
			hdmi2usbsoc_hdmi_in0_resdetection_vcounter <= (hdmi2usbsoc_hdmi_in0_resdetection_vcounter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in0_resdetection_valid_i) begin
		if (hdmi2usbsoc_hdmi_in0_resdetection_p_vsync) begin
			hdmi2usbsoc_hdmi_in0_resdetection_vcounter_st <= hdmi2usbsoc_hdmi_in0_resdetection_vcounter;
		end
	end else begin
		hdmi2usbsoc_hdmi_in0_resdetection_vcounter_st <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in0_frame_de_r <= hdmi2usbsoc_hdmi_in0_frame_de;
	hdmi2usbsoc_hdmi_in0_frame_next_de0 <= hdmi2usbsoc_hdmi_in0_frame_de;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync0 <= hdmi2usbsoc_hdmi_in0_frame_vsync;
	hdmi2usbsoc_hdmi_in0_frame_next_de1 <= hdmi2usbsoc_hdmi_in0_frame_next_de0;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync1 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync0;
	hdmi2usbsoc_hdmi_in0_frame_next_de2 <= hdmi2usbsoc_hdmi_in0_frame_next_de1;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync2 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync1;
	hdmi2usbsoc_hdmi_in0_frame_next_de3 <= hdmi2usbsoc_hdmi_in0_frame_next_de2;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync3 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync2;
	hdmi2usbsoc_hdmi_in0_frame_next_de4 <= hdmi2usbsoc_hdmi_in0_frame_next_de3;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync4 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync3;
	hdmi2usbsoc_hdmi_in0_frame_next_de5 <= hdmi2usbsoc_hdmi_in0_frame_next_de4;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync5 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync4;
	hdmi2usbsoc_hdmi_in0_frame_next_de6 <= hdmi2usbsoc_hdmi_in0_frame_next_de5;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync6 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync5;
	hdmi2usbsoc_hdmi_in0_frame_next_de7 <= hdmi2usbsoc_hdmi_in0_frame_next_de6;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync7 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync6;
	hdmi2usbsoc_hdmi_in0_frame_next_de8 <= hdmi2usbsoc_hdmi_in0_frame_next_de7;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync8 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync7;
	hdmi2usbsoc_hdmi_in0_frame_next_de9 <= hdmi2usbsoc_hdmi_in0_frame_next_de8;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync9 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync8;
	hdmi2usbsoc_hdmi_in0_frame_next_de10 <= hdmi2usbsoc_hdmi_in0_frame_next_de9;
	hdmi2usbsoc_hdmi_in0_frame_next_vsync10 <= hdmi2usbsoc_hdmi_in0_frame_next_vsync9;
	hdmi2usbsoc_hdmi_in0_frame_vsync_r <= hdmi2usbsoc_hdmi_in0_frame_next_vsync10;
	hdmi2usbsoc_hdmi_in0_frame_cur_word_valid <= 1'd0;
	if (hdmi2usbsoc_hdmi_in0_frame_new_frame) begin
		hdmi2usbsoc_hdmi_in0_frame_cur_word_valid <= (hdmi2usbsoc_hdmi_in0_frame_pack_counter == 2'd3);
		hdmi2usbsoc_hdmi_in0_frame_pack_counter <= 1'd0;
	end else begin
		if ((hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_valid & hdmi2usbsoc_hdmi_in0_frame_next_de10)) begin
			if ((hdmi2usbsoc_hdmi_in0_frame_pack_counter == 2'd3)) begin
				hdmi2usbsoc_hdmi_in0_frame_cur_word[15:0] <= hdmi2usbsoc_hdmi_in0_frame_encoded_pixel;
			end
			if ((hdmi2usbsoc_hdmi_in0_frame_pack_counter == 2'd2)) begin
				hdmi2usbsoc_hdmi_in0_frame_cur_word[31:16] <= hdmi2usbsoc_hdmi_in0_frame_encoded_pixel;
			end
			if ((hdmi2usbsoc_hdmi_in0_frame_pack_counter == 1'd1)) begin
				hdmi2usbsoc_hdmi_in0_frame_cur_word[47:32] <= hdmi2usbsoc_hdmi_in0_frame_encoded_pixel;
			end
			if ((hdmi2usbsoc_hdmi_in0_frame_pack_counter == 1'd0)) begin
				hdmi2usbsoc_hdmi_in0_frame_cur_word[63:48] <= hdmi2usbsoc_hdmi_in0_frame_encoded_pixel;
			end
			hdmi2usbsoc_hdmi_in0_frame_cur_word_valid <= (hdmi2usbsoc_hdmi_in0_frame_pack_counter == 2'd3);
			hdmi2usbsoc_hdmi_in0_frame_pack_counter <= (hdmi2usbsoc_hdmi_in0_frame_pack_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in0_frame_new_frame) begin
		hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_sof <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_frame_cur_word_valid) begin
			hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_sof <= 1'd0;
		end
	end
	if ((hdmi2usbsoc_hdmi_in0_frame_fifo_sink_valid & (~hdmi2usbsoc_hdmi_in0_frame_fifo_sink_ready))) begin
		hdmi2usbsoc_hdmi_in0_frame_pix_overflow <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_frame_pix_overflow_reset) begin
			hdmi2usbsoc_hdmi_in0_frame_pix_overflow <= 1'd0;
		end
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n0 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_valid;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n1 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n0;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n2 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n1;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n3 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n2;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n4 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n3;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n5 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n4;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n6 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n5;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n7 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n6;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n0 <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_valid & hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_first);
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n0 <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_valid & hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_last);
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n1 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n1 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n0;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n2 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n1;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n2 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n1;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n3 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n2;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n3 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n2;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n4 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n3;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n4 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n3;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n5 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n4;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n5 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n4;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n6 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n5;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n6 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n5;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n7 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n6;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n7 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n6;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_r <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_r;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_g <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_g;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_b <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_b;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_g <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_r - hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_g);
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_g <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_b - hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_sink_g);
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_ca_mult_rg <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_g * $signed({1'd0, 6'd46}));
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb_mult_bg <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_g * $signed({1'd0, 4'd15}));
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_carg_plus_cbbg <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_ca_mult_rg + hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb_mult_bg);
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_carg_plus_cbbg[24:8] + $signed({1'd0, hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_g}));
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_yraw <= ($signed({1'd0, hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_b}) - hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw);
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_yraw <= ($signed({1'd0, hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_r}) - hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw);
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r0 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cc_mult_ryraw <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_yraw * $signed({1'd0, 8'd141}));
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cd_mult_byraw <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_yraw * $signed({1'd0, 8'd166}));
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r1 <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_y <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r1 + $signed({1'd0, 5'd16}));
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cc_mult_ryraw[19:8] + $signed({1'd0, 8'd128}));
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cr <= (hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cd_mult_byraw[19:8] + $signed({1'd0, 8'd128}));
		if ((hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_y > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_y <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_y < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_y <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_y <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_y;
			end
		end
		if ((hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cb <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cb <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cb <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb;
			end
		end
		if ((hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cr > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cr <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cr < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cr <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cr <= hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cr;
			end
		end
	end
	if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n0 <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_valid;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n1 <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n0;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n2 <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n1;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n0 <= (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_valid & hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_first);
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n0 <= (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_valid & hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_last);
	end
	if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n1 <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n1 <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n0;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n2 <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n1;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n2 <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n1;
	end
	if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_ce) begin
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_y <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_y;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cb <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cb;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cr <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cr;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_y <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_y;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cb <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cr <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_y <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_y;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_cb <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_cr <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cr;
		if ((hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first | (~hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_parity))) begin
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_parity <= 1'd1;
		end else begin
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_parity <= 1'd0;
		end
		if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_parity) begin
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cb_sum <= (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cb + hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cb);
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cr_sum <= (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_sink_cr + hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cr);
		end
		if (hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_parity) begin
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_y <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_y;
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_cb_cr <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cr_mean;
		end else begin
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_y <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_y;
			hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_cb_cr <= hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cb_mean;
		end
	end
	hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_binary <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next_binary;
	hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_next;
	hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_o_r <= hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_i) begin
		hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_i <= (~hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_i);
	end
	if (hdmi_in0_pix_rst) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_d <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_data <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_raw_data1 <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_found_control <= 1'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_control_counter <= 3'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_previous_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in0_charsync0_word_sel <= 4'd0;
		hdmi2usbsoc_hdmi_in0_wer0_data_r <= 9'd0;
		hdmi2usbsoc_hdmi_in0_wer0_transition_count <= 4'd0;
		hdmi2usbsoc_hdmi_in0_wer0_is_control <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer0_is_error <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer0_period_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer0_period_done <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer0_wer_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r_updated <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_raw <= 10'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_d <= 8'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_c <= 2'd0;
		hdmi2usbsoc_hdmi_in0_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_d <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_data <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_raw_data1 <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_found_control <= 1'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_control_counter <= 3'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_previous_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in0_charsync1_word_sel <= 4'd0;
		hdmi2usbsoc_hdmi_in0_wer1_data_r <= 9'd0;
		hdmi2usbsoc_hdmi_in0_wer1_transition_count <= 4'd0;
		hdmi2usbsoc_hdmi_in0_wer1_is_control <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer1_is_error <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer1_period_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer1_period_done <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer1_wer_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r_updated <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_raw <= 10'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_d <= 8'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_c <= 2'd0;
		hdmi2usbsoc_hdmi_in0_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_d <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_data <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_raw_data1 <= 10'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_found_control <= 1'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_control_counter <= 3'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_previous_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in0_charsync2_word_sel <= 4'd0;
		hdmi2usbsoc_hdmi_in0_wer2_data_r <= 9'd0;
		hdmi2usbsoc_hdmi_in0_wer2_transition_count <= 4'd0;
		hdmi2usbsoc_hdmi_in0_wer2_is_control <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer2_is_error <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer2_period_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer2_period_done <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer2_wer_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r_updated <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_raw <= 10'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_d <= 8'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_c <= 2'd0;
		hdmi2usbsoc_hdmi_in0_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in0_chansync_chan_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_produce <= 3'd0;
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_consume <= 3'd0;
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_produce <= 3'd0;
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_consume <= 3'd0;
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_produce <= 3'd0;
		hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_consume <= 3'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_de_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_c_polarity <= 2'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_c_out <= 2'd0;
		hdmi2usbsoc_hdmi_in0_resdetection_de_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_resdetection_hcounter <= 11'd0;
		hdmi2usbsoc_hdmi_in0_resdetection_hcounter_st <= 11'd0;
		hdmi2usbsoc_hdmi_in0_resdetection_vsync_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_resdetection_vcounter <= 11'd0;
		hdmi2usbsoc_hdmi_in0_resdetection_vcounter_st <= 11'd0;
		hdmi2usbsoc_hdmi_in0_frame_de_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_y <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_source_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record0_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record1_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record2_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record3_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record4_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record5_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record6_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_record7_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_g <= 9'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_g <= 9'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_ca_mult_rg <= 17'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb_mult_bg <= 17'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_carg_plus_cbbg <= 25'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw <= 11'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_b_minus_yraw <= 12'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_r_minus_yraw <= 12'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r0 <= 11'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cc_mult_ryraw <= 20'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cd_mult_byraw <= 20'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_yraw_r1 <= 11'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_y <= 11'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cb <= 12'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_cr <= 12'sd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n3 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n4 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n5 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n6 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_valid_n7 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n3 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n3 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n4 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n4 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n5 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n5 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n6 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n6 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_first_n7 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_rgb2ycbcr_last_n7 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_y <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_source_cb_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_y <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record0_ycbcr_n_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_y <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record1_ycbcr_n_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_y <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_record2_ycbcr_n_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_parity <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cb_sum <= 9'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_cr_sum <= 9'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_valid_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_first_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_chroma_downsampler_last_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync0 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync1 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync2 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de3 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync3 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de4 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync4 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de5 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync5 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de6 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync6 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de7 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync7 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de8 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync8 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de9 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync9 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_de10 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_next_vsync10 <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_vsync_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_cur_word <= 64'd0;
		hdmi2usbsoc_hdmi_in0_frame_cur_word_valid <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_pack_counter <= 2'd0;
		hdmi2usbsoc_hdmi_in0_frame_fifo_sink_payload_sof <= 1'd0;
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q <= 10'd0;
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q_binary <= 10'd0;
		hdmi2usbsoc_hdmi_in0_frame_pix_overflow <= 1'd0;
	end
	xilinxmultiregimpl47_regs0 <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q;
	xilinxmultiregimpl47_regs1 <= xilinxmultiregimpl47_regs0;
	xilinxmultiregimpl49_regs0 <= hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_i;
	xilinxmultiregimpl49_regs1 <= xilinxmultiregimpl49_regs0;
end

always @(posedge hdmi_in0_pix2x_clk) begin
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_reset_lateness) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness <= 8'd128;
	end else begin
		if (((((~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_busy) & (~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_busy)) & (~hdmi2usbsoc_hdmi_in0_s6datacapture0_too_late)) & (~hdmi2usbsoc_hdmi_in0_s6datacapture0_too_early))) begin
			if ((hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_valid & hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_incdec)) begin
				hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness <= (hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness - 1'd1);
			end
			if ((hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_valid & (~hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_incdec))) begin
				hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness <= (hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness + 1'd1);
			end
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_pending)) begin
		if ((hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_cal | hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_ce)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_busy)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_pending)) begin
		if ((hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_cal | hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_ce)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_busy)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr <= {hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr2, hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr[9:5]};
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_i);
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_reset_lateness) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness <= 8'd128;
	end else begin
		if (((((~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_busy) & (~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_busy)) & (~hdmi2usbsoc_hdmi_in0_s6datacapture1_too_late)) & (~hdmi2usbsoc_hdmi_in0_s6datacapture1_too_early))) begin
			if ((hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_valid & hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_incdec)) begin
				hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness <= (hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness - 1'd1);
			end
			if ((hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_valid & (~hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_incdec))) begin
				hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness <= (hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness + 1'd1);
			end
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_pending)) begin
		if ((hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_cal | hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_ce)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_busy)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_pending)) begin
		if ((hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_cal | hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_ce)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_busy)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr <= {hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr2, hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr[9:5]};
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_i);
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_reset_lateness) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness <= 8'd128;
	end else begin
		if (((((~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_busy) & (~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_busy)) & (~hdmi2usbsoc_hdmi_in0_s6datacapture2_too_late)) & (~hdmi2usbsoc_hdmi_in0_s6datacapture2_too_early))) begin
			if ((hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_valid & hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_incdec)) begin
				hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness <= (hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness - 1'd1);
			end
			if ((hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_valid & (~hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_incdec))) begin
				hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness <= (hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness + 1'd1);
			end
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_pending)) begin
		if ((hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_cal | hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_ce)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_busy)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_pending)) begin
		if ((hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_cal | hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_ce)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_busy)) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr <= {hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr2, hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr[9:5]};
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_i);
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_o;
	if (hdmi_in0_pix2x_rst) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_lateness <= 8'd128;
		hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr <= 10'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_lateness <= 8'd128;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr <= 10'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_lateness <= 8'd128;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr <= 10'd0;
	end
	xilinxmultiregimpl6_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_i;
	xilinxmultiregimpl6_regs1 <= xilinxmultiregimpl6_regs0;
	xilinxmultiregimpl7_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_i;
	xilinxmultiregimpl7_regs1 <= xilinxmultiregimpl7_regs0;
	xilinxmultiregimpl8_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_i;
	xilinxmultiregimpl8_regs1 <= xilinxmultiregimpl8_regs0;
	xilinxmultiregimpl9_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_i;
	xilinxmultiregimpl9_regs1 <= xilinxmultiregimpl9_regs0;
	xilinxmultiregimpl10_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_i;
	xilinxmultiregimpl10_regs1 <= xilinxmultiregimpl10_regs0;
	xilinxmultiregimpl11_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_i;
	xilinxmultiregimpl11_regs1 <= xilinxmultiregimpl11_regs0;
	xilinxmultiregimpl13_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_i;
	xilinxmultiregimpl13_regs1 <= xilinxmultiregimpl13_regs0;
	xilinxmultiregimpl19_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_i;
	xilinxmultiregimpl19_regs1 <= xilinxmultiregimpl19_regs0;
	xilinxmultiregimpl20_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_i;
	xilinxmultiregimpl20_regs1 <= xilinxmultiregimpl20_regs0;
	xilinxmultiregimpl21_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_i;
	xilinxmultiregimpl21_regs1 <= xilinxmultiregimpl21_regs0;
	xilinxmultiregimpl22_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_i;
	xilinxmultiregimpl22_regs1 <= xilinxmultiregimpl22_regs0;
	xilinxmultiregimpl23_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_i;
	xilinxmultiregimpl23_regs1 <= xilinxmultiregimpl23_regs0;
	xilinxmultiregimpl24_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_i;
	xilinxmultiregimpl24_regs1 <= xilinxmultiregimpl24_regs0;
	xilinxmultiregimpl26_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_i;
	xilinxmultiregimpl26_regs1 <= xilinxmultiregimpl26_regs0;
	xilinxmultiregimpl32_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_i;
	xilinxmultiregimpl32_regs1 <= xilinxmultiregimpl32_regs0;
	xilinxmultiregimpl33_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_i;
	xilinxmultiregimpl33_regs1 <= xilinxmultiregimpl33_regs0;
	xilinxmultiregimpl34_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_i;
	xilinxmultiregimpl34_regs1 <= xilinxmultiregimpl34_regs0;
	xilinxmultiregimpl35_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_i;
	xilinxmultiregimpl35_regs1 <= xilinxmultiregimpl35_regs0;
	xilinxmultiregimpl36_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_i;
	xilinxmultiregimpl36_regs1 <= xilinxmultiregimpl36_regs0;
	xilinxmultiregimpl37_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_i;
	xilinxmultiregimpl37_regs1 <= xilinxmultiregimpl37_regs0;
	xilinxmultiregimpl39_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_i;
	xilinxmultiregimpl39_regs1 <= xilinxmultiregimpl39_regs0;
end

always @(posedge hdmi_in0_pix_o_clk) begin
	hdmi2usbsoc_hdmi_in0_syncpol_c0 <= hdmi2usbsoc_hdmi_in0_syncpol_data_in0_raw;
	hdmi2usbsoc_hdmi_in0_syncpol_c1 <= hdmi2usbsoc_hdmi_in0_syncpol_data_in1_raw;
	hdmi2usbsoc_hdmi_in0_syncpol_c2 <= hdmi2usbsoc_hdmi_in0_syncpol_data_in2_raw;
	if (hdmi_in0_pix_o_rst) begin
		hdmi2usbsoc_hdmi_in0_syncpol_c0 <= 10'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_c1 <= 10'd0;
		hdmi2usbsoc_hdmi_in0_syncpol_c2 <= 10'd0;
	end
end

always @(posedge hdmi_in1_pix_clk) begin
	hdmi2usbsoc_hdmi_in1_s6datacapture0_d <= hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr;
	hdmi2usbsoc_hdmi_in1_charsync0_raw_data1 <= hdmi2usbsoc_hdmi_in1_charsync0_raw_data;
	hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd0;
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[9:0] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[9:0] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[9:0] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[9:0] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 1'd0;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[10:1] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[10:1] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[10:1] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[10:1] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 1'd1;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[11:2] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[11:2] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[11:2] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[11:2] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 2'd2;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[12:3] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[12:3] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[12:3] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[12:3] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 2'd3;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[13:4] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[13:4] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[13:4] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[13:4] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 3'd4;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[14:5] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[14:5] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[14:5] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[14:5] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 3'd5;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[15:6] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[15:6] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[15:6] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[15:6] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 3'd6;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[16:7] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[16:7] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[16:7] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[16:7] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 3'd7;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[17:8] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[17:8] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[17:8] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[17:8] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 4'd8;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync0_raw[18:9] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[18:9] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[18:9] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync0_raw[18:9] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 4'd9;
	end
	if ((hdmi2usbsoc_hdmi_in1_charsync0_found_control & (hdmi2usbsoc_hdmi_in1_charsync0_control_position == hdmi2usbsoc_hdmi_in1_charsync0_previous_control_position))) begin
		if ((hdmi2usbsoc_hdmi_in1_charsync0_control_counter == 3'd7)) begin
			hdmi2usbsoc_hdmi_in1_charsync0_control_counter <= 1'd0;
			hdmi2usbsoc_hdmi_in1_charsync0_synced <= 1'd1;
			hdmi2usbsoc_hdmi_in1_charsync0_word_sel <= hdmi2usbsoc_hdmi_in1_charsync0_control_position;
		end else begin
			hdmi2usbsoc_hdmi_in1_charsync0_control_counter <= (hdmi2usbsoc_hdmi_in1_charsync0_control_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_in1_charsync0_control_counter <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in1_charsync0_previous_control_position <= hdmi2usbsoc_hdmi_in1_charsync0_control_position;
	hdmi2usbsoc_hdmi_in1_charsync0_data <= (hdmi2usbsoc_hdmi_in1_charsync0_raw >>> hdmi2usbsoc_hdmi_in1_charsync0_word_sel);
	hdmi2usbsoc_hdmi_in1_wer0_data_r <= hdmi2usbsoc_hdmi_in1_wer0_data[8:0];
	hdmi2usbsoc_hdmi_in1_wer0_transition_count <= (((((((hdmi2usbsoc_hdmi_in1_wer0_transitions[0] + hdmi2usbsoc_hdmi_in1_wer0_transitions[1]) + hdmi2usbsoc_hdmi_in1_wer0_transitions[2]) + hdmi2usbsoc_hdmi_in1_wer0_transitions[3]) + hdmi2usbsoc_hdmi_in1_wer0_transitions[4]) + hdmi2usbsoc_hdmi_in1_wer0_transitions[5]) + hdmi2usbsoc_hdmi_in1_wer0_transitions[6]) + hdmi2usbsoc_hdmi_in1_wer0_transitions[7]);
	hdmi2usbsoc_hdmi_in1_wer0_is_control <= ((((hdmi2usbsoc_hdmi_in1_wer0_data_r == 10'd852) | (hdmi2usbsoc_hdmi_in1_wer0_data_r == 8'd171)) | (hdmi2usbsoc_hdmi_in1_wer0_data_r == 9'd340)) | (hdmi2usbsoc_hdmi_in1_wer0_data_r == 10'd683));
	hdmi2usbsoc_hdmi_in1_wer0_is_error <= ((hdmi2usbsoc_hdmi_in1_wer0_transition_count > 3'd4) & (~hdmi2usbsoc_hdmi_in1_wer0_is_control));
	{hdmi2usbsoc_hdmi_in1_wer0_period_done, hdmi2usbsoc_hdmi_in1_wer0_period_counter} <= (hdmi2usbsoc_hdmi_in1_wer0_period_counter + 1'd1);
	hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r_updated <= hdmi2usbsoc_hdmi_in1_wer0_period_done;
	if (hdmi2usbsoc_hdmi_in1_wer0_period_done) begin
		hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r <= hdmi2usbsoc_hdmi_in1_wer0_wer_counter;
		hdmi2usbsoc_hdmi_in1_wer0_wer_counter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_wer0_is_error) begin
			hdmi2usbsoc_hdmi_in1_wer0_wer_counter <= (hdmi2usbsoc_hdmi_in1_wer0_wer_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in1_wer0_i) begin
		hdmi2usbsoc_hdmi_in1_wer0_toggle_i <= (~hdmi2usbsoc_hdmi_in1_wer0_toggle_i);
	end
	hdmi2usbsoc_hdmi_in1_decoding0_output_de <= 1'd1;
	if ((hdmi2usbsoc_hdmi_in1_decoding0_input == 10'd852)) begin
		hdmi2usbsoc_hdmi_in1_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_c <= 1'd0;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding0_input == 8'd171)) begin
		hdmi2usbsoc_hdmi_in1_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_c <= 1'd1;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding0_input == 9'd340)) begin
		hdmi2usbsoc_hdmi_in1_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_c <= 2'd2;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding0_input == 10'd683)) begin
		hdmi2usbsoc_hdmi_in1_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_c <= 2'd3;
	end
	hdmi2usbsoc_hdmi_in1_decoding0_output_raw <= hdmi2usbsoc_hdmi_in1_decoding0_input;
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[0] <= (hdmi2usbsoc_hdmi_in1_decoding0_input[0] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[9]);
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[1] <= ((hdmi2usbsoc_hdmi_in1_decoding0_input[1] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[0]) ^ (~hdmi2usbsoc_hdmi_in1_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[2] <= ((hdmi2usbsoc_hdmi_in1_decoding0_input[2] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[1]) ^ (~hdmi2usbsoc_hdmi_in1_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[3] <= ((hdmi2usbsoc_hdmi_in1_decoding0_input[3] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[2]) ^ (~hdmi2usbsoc_hdmi_in1_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[4] <= ((hdmi2usbsoc_hdmi_in1_decoding0_input[4] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[3]) ^ (~hdmi2usbsoc_hdmi_in1_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[5] <= ((hdmi2usbsoc_hdmi_in1_decoding0_input[5] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[4]) ^ (~hdmi2usbsoc_hdmi_in1_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[6] <= ((hdmi2usbsoc_hdmi_in1_decoding0_input[6] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[5]) ^ (~hdmi2usbsoc_hdmi_in1_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding0_output_d[7] <= ((hdmi2usbsoc_hdmi_in1_decoding0_input[7] ^ hdmi2usbsoc_hdmi_in1_decoding0_input[6]) ^ (~hdmi2usbsoc_hdmi_in1_decoding0_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding0_valid_o <= hdmi2usbsoc_hdmi_in1_decoding0_valid_i;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_d <= hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr;
	hdmi2usbsoc_hdmi_in1_charsync1_raw_data1 <= hdmi2usbsoc_hdmi_in1_charsync1_raw_data;
	hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd0;
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[9:0] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[9:0] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[9:0] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[9:0] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 1'd0;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[10:1] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[10:1] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[10:1] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[10:1] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 1'd1;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[11:2] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[11:2] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[11:2] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[11:2] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 2'd2;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[12:3] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[12:3] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[12:3] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[12:3] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 2'd3;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[13:4] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[13:4] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[13:4] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[13:4] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 3'd4;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[14:5] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[14:5] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[14:5] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[14:5] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 3'd5;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[15:6] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[15:6] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[15:6] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[15:6] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 3'd6;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[16:7] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[16:7] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[16:7] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[16:7] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 3'd7;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[17:8] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[17:8] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[17:8] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[17:8] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 4'd8;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync1_raw[18:9] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[18:9] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[18:9] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync1_raw[18:9] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 4'd9;
	end
	if ((hdmi2usbsoc_hdmi_in1_charsync1_found_control & (hdmi2usbsoc_hdmi_in1_charsync1_control_position == hdmi2usbsoc_hdmi_in1_charsync1_previous_control_position))) begin
		if ((hdmi2usbsoc_hdmi_in1_charsync1_control_counter == 3'd7)) begin
			hdmi2usbsoc_hdmi_in1_charsync1_control_counter <= 1'd0;
			hdmi2usbsoc_hdmi_in1_charsync1_synced <= 1'd1;
			hdmi2usbsoc_hdmi_in1_charsync1_word_sel <= hdmi2usbsoc_hdmi_in1_charsync1_control_position;
		end else begin
			hdmi2usbsoc_hdmi_in1_charsync1_control_counter <= (hdmi2usbsoc_hdmi_in1_charsync1_control_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_in1_charsync1_control_counter <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in1_charsync1_previous_control_position <= hdmi2usbsoc_hdmi_in1_charsync1_control_position;
	hdmi2usbsoc_hdmi_in1_charsync1_data <= (hdmi2usbsoc_hdmi_in1_charsync1_raw >>> hdmi2usbsoc_hdmi_in1_charsync1_word_sel);
	hdmi2usbsoc_hdmi_in1_wer1_data_r <= hdmi2usbsoc_hdmi_in1_wer1_data[8:0];
	hdmi2usbsoc_hdmi_in1_wer1_transition_count <= (((((((hdmi2usbsoc_hdmi_in1_wer1_transitions[0] + hdmi2usbsoc_hdmi_in1_wer1_transitions[1]) + hdmi2usbsoc_hdmi_in1_wer1_transitions[2]) + hdmi2usbsoc_hdmi_in1_wer1_transitions[3]) + hdmi2usbsoc_hdmi_in1_wer1_transitions[4]) + hdmi2usbsoc_hdmi_in1_wer1_transitions[5]) + hdmi2usbsoc_hdmi_in1_wer1_transitions[6]) + hdmi2usbsoc_hdmi_in1_wer1_transitions[7]);
	hdmi2usbsoc_hdmi_in1_wer1_is_control <= ((((hdmi2usbsoc_hdmi_in1_wer1_data_r == 10'd852) | (hdmi2usbsoc_hdmi_in1_wer1_data_r == 8'd171)) | (hdmi2usbsoc_hdmi_in1_wer1_data_r == 9'd340)) | (hdmi2usbsoc_hdmi_in1_wer1_data_r == 10'd683));
	hdmi2usbsoc_hdmi_in1_wer1_is_error <= ((hdmi2usbsoc_hdmi_in1_wer1_transition_count > 3'd4) & (~hdmi2usbsoc_hdmi_in1_wer1_is_control));
	{hdmi2usbsoc_hdmi_in1_wer1_period_done, hdmi2usbsoc_hdmi_in1_wer1_period_counter} <= (hdmi2usbsoc_hdmi_in1_wer1_period_counter + 1'd1);
	hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r_updated <= hdmi2usbsoc_hdmi_in1_wer1_period_done;
	if (hdmi2usbsoc_hdmi_in1_wer1_period_done) begin
		hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r <= hdmi2usbsoc_hdmi_in1_wer1_wer_counter;
		hdmi2usbsoc_hdmi_in1_wer1_wer_counter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_wer1_is_error) begin
			hdmi2usbsoc_hdmi_in1_wer1_wer_counter <= (hdmi2usbsoc_hdmi_in1_wer1_wer_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in1_wer1_i) begin
		hdmi2usbsoc_hdmi_in1_wer1_toggle_i <= (~hdmi2usbsoc_hdmi_in1_wer1_toggle_i);
	end
	hdmi2usbsoc_hdmi_in1_decoding1_output_de <= 1'd1;
	if ((hdmi2usbsoc_hdmi_in1_decoding1_input == 10'd852)) begin
		hdmi2usbsoc_hdmi_in1_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_c <= 1'd0;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding1_input == 8'd171)) begin
		hdmi2usbsoc_hdmi_in1_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_c <= 1'd1;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding1_input == 9'd340)) begin
		hdmi2usbsoc_hdmi_in1_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_c <= 2'd2;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding1_input == 10'd683)) begin
		hdmi2usbsoc_hdmi_in1_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_c <= 2'd3;
	end
	hdmi2usbsoc_hdmi_in1_decoding1_output_raw <= hdmi2usbsoc_hdmi_in1_decoding1_input;
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[0] <= (hdmi2usbsoc_hdmi_in1_decoding1_input[0] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[9]);
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[1] <= ((hdmi2usbsoc_hdmi_in1_decoding1_input[1] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[0]) ^ (~hdmi2usbsoc_hdmi_in1_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[2] <= ((hdmi2usbsoc_hdmi_in1_decoding1_input[2] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[1]) ^ (~hdmi2usbsoc_hdmi_in1_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[3] <= ((hdmi2usbsoc_hdmi_in1_decoding1_input[3] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[2]) ^ (~hdmi2usbsoc_hdmi_in1_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[4] <= ((hdmi2usbsoc_hdmi_in1_decoding1_input[4] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[3]) ^ (~hdmi2usbsoc_hdmi_in1_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[5] <= ((hdmi2usbsoc_hdmi_in1_decoding1_input[5] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[4]) ^ (~hdmi2usbsoc_hdmi_in1_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[6] <= ((hdmi2usbsoc_hdmi_in1_decoding1_input[6] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[5]) ^ (~hdmi2usbsoc_hdmi_in1_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding1_output_d[7] <= ((hdmi2usbsoc_hdmi_in1_decoding1_input[7] ^ hdmi2usbsoc_hdmi_in1_decoding1_input[6]) ^ (~hdmi2usbsoc_hdmi_in1_decoding1_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding1_valid_o <= hdmi2usbsoc_hdmi_in1_decoding1_valid_i;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_d <= hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr;
	hdmi2usbsoc_hdmi_in1_charsync2_raw_data1 <= hdmi2usbsoc_hdmi_in1_charsync2_raw_data;
	hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd0;
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[9:0] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[9:0] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[9:0] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[9:0] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 1'd0;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[10:1] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[10:1] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[10:1] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[10:1] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 1'd1;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[11:2] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[11:2] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[11:2] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[11:2] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 2'd2;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[12:3] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[12:3] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[12:3] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[12:3] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 2'd3;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[13:4] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[13:4] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[13:4] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[13:4] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 3'd4;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[14:5] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[14:5] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[14:5] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[14:5] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 3'd5;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[15:6] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[15:6] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[15:6] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[15:6] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 3'd6;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[16:7] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[16:7] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[16:7] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[16:7] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 3'd7;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[17:8] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[17:8] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[17:8] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[17:8] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 4'd8;
	end
	if (((((hdmi2usbsoc_hdmi_in1_charsync2_raw[18:9] == 10'd852) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[18:9] == 8'd171)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[18:9] == 9'd340)) | (hdmi2usbsoc_hdmi_in1_charsync2_raw[18:9] == 10'd683))) begin
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd1;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 4'd9;
	end
	if ((hdmi2usbsoc_hdmi_in1_charsync2_found_control & (hdmi2usbsoc_hdmi_in1_charsync2_control_position == hdmi2usbsoc_hdmi_in1_charsync2_previous_control_position))) begin
		if ((hdmi2usbsoc_hdmi_in1_charsync2_control_counter == 3'd7)) begin
			hdmi2usbsoc_hdmi_in1_charsync2_control_counter <= 1'd0;
			hdmi2usbsoc_hdmi_in1_charsync2_synced <= 1'd1;
			hdmi2usbsoc_hdmi_in1_charsync2_word_sel <= hdmi2usbsoc_hdmi_in1_charsync2_control_position;
		end else begin
			hdmi2usbsoc_hdmi_in1_charsync2_control_counter <= (hdmi2usbsoc_hdmi_in1_charsync2_control_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_in1_charsync2_control_counter <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in1_charsync2_previous_control_position <= hdmi2usbsoc_hdmi_in1_charsync2_control_position;
	hdmi2usbsoc_hdmi_in1_charsync2_data <= (hdmi2usbsoc_hdmi_in1_charsync2_raw >>> hdmi2usbsoc_hdmi_in1_charsync2_word_sel);
	hdmi2usbsoc_hdmi_in1_wer2_data_r <= hdmi2usbsoc_hdmi_in1_wer2_data[8:0];
	hdmi2usbsoc_hdmi_in1_wer2_transition_count <= (((((((hdmi2usbsoc_hdmi_in1_wer2_transitions[0] + hdmi2usbsoc_hdmi_in1_wer2_transitions[1]) + hdmi2usbsoc_hdmi_in1_wer2_transitions[2]) + hdmi2usbsoc_hdmi_in1_wer2_transitions[3]) + hdmi2usbsoc_hdmi_in1_wer2_transitions[4]) + hdmi2usbsoc_hdmi_in1_wer2_transitions[5]) + hdmi2usbsoc_hdmi_in1_wer2_transitions[6]) + hdmi2usbsoc_hdmi_in1_wer2_transitions[7]);
	hdmi2usbsoc_hdmi_in1_wer2_is_control <= ((((hdmi2usbsoc_hdmi_in1_wer2_data_r == 10'd852) | (hdmi2usbsoc_hdmi_in1_wer2_data_r == 8'd171)) | (hdmi2usbsoc_hdmi_in1_wer2_data_r == 9'd340)) | (hdmi2usbsoc_hdmi_in1_wer2_data_r == 10'd683));
	hdmi2usbsoc_hdmi_in1_wer2_is_error <= ((hdmi2usbsoc_hdmi_in1_wer2_transition_count > 3'd4) & (~hdmi2usbsoc_hdmi_in1_wer2_is_control));
	{hdmi2usbsoc_hdmi_in1_wer2_period_done, hdmi2usbsoc_hdmi_in1_wer2_period_counter} <= (hdmi2usbsoc_hdmi_in1_wer2_period_counter + 1'd1);
	hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r_updated <= hdmi2usbsoc_hdmi_in1_wer2_period_done;
	if (hdmi2usbsoc_hdmi_in1_wer2_period_done) begin
		hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r <= hdmi2usbsoc_hdmi_in1_wer2_wer_counter;
		hdmi2usbsoc_hdmi_in1_wer2_wer_counter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_wer2_is_error) begin
			hdmi2usbsoc_hdmi_in1_wer2_wer_counter <= (hdmi2usbsoc_hdmi_in1_wer2_wer_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in1_wer2_i) begin
		hdmi2usbsoc_hdmi_in1_wer2_toggle_i <= (~hdmi2usbsoc_hdmi_in1_wer2_toggle_i);
	end
	hdmi2usbsoc_hdmi_in1_decoding2_output_de <= 1'd1;
	if ((hdmi2usbsoc_hdmi_in1_decoding2_input == 10'd852)) begin
		hdmi2usbsoc_hdmi_in1_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_c <= 1'd0;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding2_input == 8'd171)) begin
		hdmi2usbsoc_hdmi_in1_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_c <= 1'd1;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding2_input == 9'd340)) begin
		hdmi2usbsoc_hdmi_in1_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_c <= 2'd2;
	end
	if ((hdmi2usbsoc_hdmi_in1_decoding2_input == 10'd683)) begin
		hdmi2usbsoc_hdmi_in1_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_c <= 2'd3;
	end
	hdmi2usbsoc_hdmi_in1_decoding2_output_raw <= hdmi2usbsoc_hdmi_in1_decoding2_input;
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[0] <= (hdmi2usbsoc_hdmi_in1_decoding2_input[0] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[9]);
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[1] <= ((hdmi2usbsoc_hdmi_in1_decoding2_input[1] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[0]) ^ (~hdmi2usbsoc_hdmi_in1_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[2] <= ((hdmi2usbsoc_hdmi_in1_decoding2_input[2] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[1]) ^ (~hdmi2usbsoc_hdmi_in1_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[3] <= ((hdmi2usbsoc_hdmi_in1_decoding2_input[3] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[2]) ^ (~hdmi2usbsoc_hdmi_in1_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[4] <= ((hdmi2usbsoc_hdmi_in1_decoding2_input[4] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[3]) ^ (~hdmi2usbsoc_hdmi_in1_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[5] <= ((hdmi2usbsoc_hdmi_in1_decoding2_input[5] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[4]) ^ (~hdmi2usbsoc_hdmi_in1_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[6] <= ((hdmi2usbsoc_hdmi_in1_decoding2_input[6] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[5]) ^ (~hdmi2usbsoc_hdmi_in1_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding2_output_d[7] <= ((hdmi2usbsoc_hdmi_in1_decoding2_input[7] ^ hdmi2usbsoc_hdmi_in1_decoding2_input[6]) ^ (~hdmi2usbsoc_hdmi_in1_decoding2_input[8]));
	hdmi2usbsoc_hdmi_in1_decoding2_valid_o <= hdmi2usbsoc_hdmi_in1_decoding2_valid_i;
	if ((~hdmi2usbsoc_hdmi_in1_chansync_valid_i)) begin
		hdmi2usbsoc_hdmi_in1_chansync_chan_synced <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_chansync_some_control) begin
			if (hdmi2usbsoc_hdmi_in1_chansync_all_control) begin
				hdmi2usbsoc_hdmi_in1_chansync_chan_synced <= 1'd1;
			end else begin
				hdmi2usbsoc_hdmi_in1_chansync_chan_synced <= 1'd0;
			end
		end
	end
	hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_produce <= (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_produce + 1'd1);
	if (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_re) begin
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_consume <= (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_consume + 1'd1);
	end
	hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_produce <= (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_produce + 1'd1);
	if (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_re) begin
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_consume <= (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_consume + 1'd1);
	end
	hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_produce <= (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_produce + 1'd1);
	if (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_re) begin
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_consume <= (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_consume + 1'd1);
	end
	hdmi2usbsoc_hdmi_in1_syncpol_valid_o <= hdmi2usbsoc_hdmi_in1_syncpol_valid_i;
	hdmi2usbsoc_hdmi_in1_syncpol_r <= hdmi2usbsoc_hdmi_in1_syncpol_data_in2_d;
	hdmi2usbsoc_hdmi_in1_syncpol_g <= hdmi2usbsoc_hdmi_in1_syncpol_data_in1_d;
	hdmi2usbsoc_hdmi_in1_syncpol_b <= hdmi2usbsoc_hdmi_in1_syncpol_data_in0_d;
	hdmi2usbsoc_hdmi_in1_syncpol_de_r <= hdmi2usbsoc_hdmi_in1_syncpol_data_in0_de;
	if ((hdmi2usbsoc_hdmi_in1_syncpol_de_r & (~hdmi2usbsoc_hdmi_in1_syncpol_data_in0_de))) begin
		hdmi2usbsoc_hdmi_in1_syncpol_c_polarity <= hdmi2usbsoc_hdmi_in1_syncpol_data_in0_c;
		hdmi2usbsoc_hdmi_in1_syncpol_c_out <= 1'd0;
	end else begin
		hdmi2usbsoc_hdmi_in1_syncpol_c_out <= (hdmi2usbsoc_hdmi_in1_syncpol_data_in0_c ^ hdmi2usbsoc_hdmi_in1_syncpol_c_polarity);
	end
	hdmi2usbsoc_hdmi_in1_resdetection_de_r <= hdmi2usbsoc_hdmi_in1_resdetection_de;
	if ((hdmi2usbsoc_hdmi_in1_resdetection_valid_i & hdmi2usbsoc_hdmi_in1_resdetection_de)) begin
		hdmi2usbsoc_hdmi_in1_resdetection_hcounter <= (hdmi2usbsoc_hdmi_in1_resdetection_hcounter + 1'd1);
	end else begin
		hdmi2usbsoc_hdmi_in1_resdetection_hcounter <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_in1_resdetection_valid_i) begin
		if (hdmi2usbsoc_hdmi_in1_resdetection_pn_de) begin
			hdmi2usbsoc_hdmi_in1_resdetection_hcounter_st <= hdmi2usbsoc_hdmi_in1_resdetection_hcounter;
		end
	end else begin
		hdmi2usbsoc_hdmi_in1_resdetection_hcounter_st <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in1_resdetection_vsync_r <= hdmi2usbsoc_hdmi_in1_resdetection_vsync;
	if ((hdmi2usbsoc_hdmi_in1_resdetection_valid_i & hdmi2usbsoc_hdmi_in1_resdetection_p_vsync)) begin
		hdmi2usbsoc_hdmi_in1_resdetection_vcounter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_resdetection_pn_de) begin
			hdmi2usbsoc_hdmi_in1_resdetection_vcounter <= (hdmi2usbsoc_hdmi_in1_resdetection_vcounter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in1_resdetection_valid_i) begin
		if (hdmi2usbsoc_hdmi_in1_resdetection_p_vsync) begin
			hdmi2usbsoc_hdmi_in1_resdetection_vcounter_st <= hdmi2usbsoc_hdmi_in1_resdetection_vcounter;
		end
	end else begin
		hdmi2usbsoc_hdmi_in1_resdetection_vcounter_st <= 1'd0;
	end
	hdmi2usbsoc_hdmi_in1_frame_de_r <= hdmi2usbsoc_hdmi_in1_frame_de;
	hdmi2usbsoc_hdmi_in1_frame_next_de0 <= hdmi2usbsoc_hdmi_in1_frame_de;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync0 <= hdmi2usbsoc_hdmi_in1_frame_vsync;
	hdmi2usbsoc_hdmi_in1_frame_next_de1 <= hdmi2usbsoc_hdmi_in1_frame_next_de0;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync1 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync0;
	hdmi2usbsoc_hdmi_in1_frame_next_de2 <= hdmi2usbsoc_hdmi_in1_frame_next_de1;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync2 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync1;
	hdmi2usbsoc_hdmi_in1_frame_next_de3 <= hdmi2usbsoc_hdmi_in1_frame_next_de2;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync3 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync2;
	hdmi2usbsoc_hdmi_in1_frame_next_de4 <= hdmi2usbsoc_hdmi_in1_frame_next_de3;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync4 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync3;
	hdmi2usbsoc_hdmi_in1_frame_next_de5 <= hdmi2usbsoc_hdmi_in1_frame_next_de4;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync5 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync4;
	hdmi2usbsoc_hdmi_in1_frame_next_de6 <= hdmi2usbsoc_hdmi_in1_frame_next_de5;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync6 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync5;
	hdmi2usbsoc_hdmi_in1_frame_next_de7 <= hdmi2usbsoc_hdmi_in1_frame_next_de6;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync7 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync6;
	hdmi2usbsoc_hdmi_in1_frame_next_de8 <= hdmi2usbsoc_hdmi_in1_frame_next_de7;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync8 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync7;
	hdmi2usbsoc_hdmi_in1_frame_next_de9 <= hdmi2usbsoc_hdmi_in1_frame_next_de8;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync9 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync8;
	hdmi2usbsoc_hdmi_in1_frame_next_de10 <= hdmi2usbsoc_hdmi_in1_frame_next_de9;
	hdmi2usbsoc_hdmi_in1_frame_next_vsync10 <= hdmi2usbsoc_hdmi_in1_frame_next_vsync9;
	hdmi2usbsoc_hdmi_in1_frame_vsync_r <= hdmi2usbsoc_hdmi_in1_frame_next_vsync10;
	hdmi2usbsoc_hdmi_in1_frame_cur_word_valid <= 1'd0;
	if (hdmi2usbsoc_hdmi_in1_frame_new_frame) begin
		hdmi2usbsoc_hdmi_in1_frame_cur_word_valid <= (hdmi2usbsoc_hdmi_in1_frame_pack_counter == 2'd3);
		hdmi2usbsoc_hdmi_in1_frame_pack_counter <= 1'd0;
	end else begin
		if ((hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_valid & hdmi2usbsoc_hdmi_in1_frame_next_de10)) begin
			if ((hdmi2usbsoc_hdmi_in1_frame_pack_counter == 2'd3)) begin
				hdmi2usbsoc_hdmi_in1_frame_cur_word[15:0] <= hdmi2usbsoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((hdmi2usbsoc_hdmi_in1_frame_pack_counter == 2'd2)) begin
				hdmi2usbsoc_hdmi_in1_frame_cur_word[31:16] <= hdmi2usbsoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((hdmi2usbsoc_hdmi_in1_frame_pack_counter == 1'd1)) begin
				hdmi2usbsoc_hdmi_in1_frame_cur_word[47:32] <= hdmi2usbsoc_hdmi_in1_frame_encoded_pixel;
			end
			if ((hdmi2usbsoc_hdmi_in1_frame_pack_counter == 1'd0)) begin
				hdmi2usbsoc_hdmi_in1_frame_cur_word[63:48] <= hdmi2usbsoc_hdmi_in1_frame_encoded_pixel;
			end
			hdmi2usbsoc_hdmi_in1_frame_cur_word_valid <= (hdmi2usbsoc_hdmi_in1_frame_pack_counter == 2'd3);
			hdmi2usbsoc_hdmi_in1_frame_pack_counter <= (hdmi2usbsoc_hdmi_in1_frame_pack_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in1_frame_new_frame) begin
		hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_sof <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_frame_cur_word_valid) begin
			hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_sof <= 1'd0;
		end
	end
	if ((hdmi2usbsoc_hdmi_in1_frame_fifo_sink_valid & (~hdmi2usbsoc_hdmi_in1_frame_fifo_sink_ready))) begin
		hdmi2usbsoc_hdmi_in1_frame_pix_overflow <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_frame_pix_overflow_reset) begin
			hdmi2usbsoc_hdmi_in1_frame_pix_overflow <= 1'd0;
		end
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n0 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_valid;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n1 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n0;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n2 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n1;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n3 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n2;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n4 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n3;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n5 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n4;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n6 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n5;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n7 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n6;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n0 <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_valid & hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_first);
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n0 <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_valid & hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_last);
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n1 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n1 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n0;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n2 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n1;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n2 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n1;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n3 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n2;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n3 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n2;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n4 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n3;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n4 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n3;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n5 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n4;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n5 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n4;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n6 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n5;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n6 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n5;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n7 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n6;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n7 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n6;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_r <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_r;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_g <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_g;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_b <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_b;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_g <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_r - hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_g);
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_g <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_b - hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_sink_g);
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_ca_mult_rg <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_g * $signed({1'd0, 6'd46}));
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb_mult_bg <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_g * $signed({1'd0, 4'd15}));
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_carg_plus_cbbg <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_ca_mult_rg + hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb_mult_bg);
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_carg_plus_cbbg[24:8] + $signed({1'd0, hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_g}));
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_yraw <= ($signed({1'd0, hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_b}) - hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw);
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_yraw <= ($signed({1'd0, hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_r}) - hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw);
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r0 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cc_mult_ryraw <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_yraw * $signed({1'd0, 8'd141}));
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cd_mult_byraw <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_yraw * $signed({1'd0, 8'd166}));
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r1 <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_y <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r1 + $signed({1'd0, 5'd16}));
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cc_mult_ryraw[19:8] + $signed({1'd0, 8'd128}));
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cr <= (hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cd_mult_byraw[19:8] + $signed({1'd0, 8'd128}));
		if ((hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_y > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_y <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_y < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_y <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_y <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_y;
			end
		end
		if ((hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cb <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cb <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cb <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb;
			end
		end
		if ((hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cr > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cr <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cr < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cr <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cr <= hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cr;
			end
		end
	end
	if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n0 <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_valid;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n1 <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n0;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n2 <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n1;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n0 <= (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_valid & hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_first);
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n0 <= (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_valid & hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_last);
	end
	if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n1 <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n1 <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n0;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_pipe_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n2 <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n1;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n2 <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n1;
	end
	if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_ce) begin
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_y <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_y;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cb <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cb;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cr <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cr;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_y <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_y;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cb <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cr <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_y <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_y;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_cb <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_cr <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cr;
		if ((hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first | (~hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_parity))) begin
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_parity <= 1'd1;
		end else begin
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_parity <= 1'd0;
		end
		if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_parity) begin
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cb_sum <= (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cb + hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cb);
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cr_sum <= (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_sink_cr + hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cr);
		end
		if (hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_parity) begin
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_y <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_y;
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_cb_cr <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cr_mean;
		end else begin
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_y <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_y;
			hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_cb_cr <= hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cb_mean;
		end
	end
	hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_binary <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next_binary;
	hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_next;
	hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_o_r <= hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_i) begin
		hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_i <= (~hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_i);
	end
	if (hdmi_in1_pix_rst) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_d <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_data <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_raw_data1 <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_found_control <= 1'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_control_counter <= 3'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_previous_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in1_charsync0_word_sel <= 4'd0;
		hdmi2usbsoc_hdmi_in1_wer0_data_r <= 9'd0;
		hdmi2usbsoc_hdmi_in1_wer0_transition_count <= 4'd0;
		hdmi2usbsoc_hdmi_in1_wer0_is_control <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer0_is_error <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer0_period_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer0_period_done <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer0_wer_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r_updated <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_raw <= 10'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_d <= 8'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_c <= 2'd0;
		hdmi2usbsoc_hdmi_in1_decoding0_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_d <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_data <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_raw_data1 <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_found_control <= 1'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_control_counter <= 3'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_previous_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in1_charsync1_word_sel <= 4'd0;
		hdmi2usbsoc_hdmi_in1_wer1_data_r <= 9'd0;
		hdmi2usbsoc_hdmi_in1_wer1_transition_count <= 4'd0;
		hdmi2usbsoc_hdmi_in1_wer1_is_control <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer1_is_error <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer1_period_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer1_period_done <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer1_wer_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r_updated <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_raw <= 10'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_d <= 8'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_c <= 2'd0;
		hdmi2usbsoc_hdmi_in1_decoding1_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_d <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_data <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_raw_data1 <= 10'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_found_control <= 1'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_control_counter <= 3'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_previous_control_position <= 4'd0;
		hdmi2usbsoc_hdmi_in1_charsync2_word_sel <= 4'd0;
		hdmi2usbsoc_hdmi_in1_wer2_data_r <= 9'd0;
		hdmi2usbsoc_hdmi_in1_wer2_transition_count <= 4'd0;
		hdmi2usbsoc_hdmi_in1_wer2_is_control <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer2_is_error <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer2_period_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer2_period_done <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer2_wer_counter <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r_updated <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_raw <= 10'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_d <= 8'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_c <= 2'd0;
		hdmi2usbsoc_hdmi_in1_decoding2_output_de <= 1'd0;
		hdmi2usbsoc_hdmi_in1_chansync_chan_synced <= 1'd0;
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_produce <= 3'd0;
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_consume <= 3'd0;
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_produce <= 3'd0;
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_consume <= 3'd0;
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_produce <= 3'd0;
		hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_consume <= 3'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_valid_o <= 1'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_de_r <= 1'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_c_polarity <= 2'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_c_out <= 2'd0;
		hdmi2usbsoc_hdmi_in1_resdetection_de_r <= 1'd0;
		hdmi2usbsoc_hdmi_in1_resdetection_hcounter <= 11'd0;
		hdmi2usbsoc_hdmi_in1_resdetection_hcounter_st <= 11'd0;
		hdmi2usbsoc_hdmi_in1_resdetection_vsync_r <= 1'd0;
		hdmi2usbsoc_hdmi_in1_resdetection_vcounter <= 11'd0;
		hdmi2usbsoc_hdmi_in1_resdetection_vcounter_st <= 11'd0;
		hdmi2usbsoc_hdmi_in1_frame_de_r <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_y <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_source_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record0_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record1_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record2_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record3_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record4_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record5_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record6_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_r <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_g <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_record7_rgb_n_b <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_g <= 9'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_g <= 9'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_ca_mult_rg <= 17'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb_mult_bg <= 17'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_carg_plus_cbbg <= 25'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw <= 11'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_b_minus_yraw <= 12'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_r_minus_yraw <= 12'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r0 <= 11'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cc_mult_ryraw <= 20'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cd_mult_byraw <= 20'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_yraw_r1 <= 11'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_y <= 11'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cb <= 12'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_cr <= 12'sd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n3 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n4 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n5 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n6 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_valid_n7 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n3 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n3 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n4 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n4 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n5 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n5 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n6 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n6 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_first_n7 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_rgb2ycbcr_last_n7 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_y <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_source_cb_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_y <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record0_ycbcr_n_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_y <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record1_ycbcr_n_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_y <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_cb <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_record2_ycbcr_n_cr <= 8'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_parity <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cb_sum <= 9'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_cr_sum <= 9'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_valid_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_first_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_chroma_downsampler_last_n2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync0 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync1 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync2 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de3 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync3 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de4 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync4 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de5 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync5 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de6 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync6 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de7 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync7 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de8 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync8 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de9 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync9 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_de10 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_next_vsync10 <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_vsync_r <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_cur_word <= 64'd0;
		hdmi2usbsoc_hdmi_in1_frame_cur_word_valid <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_pack_counter <= 2'd0;
		hdmi2usbsoc_hdmi_in1_frame_fifo_sink_payload_sof <= 1'd0;
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q <= 10'd0;
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q_binary <= 10'd0;
		hdmi2usbsoc_hdmi_in1_frame_pix_overflow <= 1'd0;
	end
	xilinxmultiregimpl97_regs0 <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q;
	xilinxmultiregimpl97_regs1 <= xilinxmultiregimpl97_regs0;
	xilinxmultiregimpl99_regs0 <= hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_i;
	xilinxmultiregimpl99_regs1 <= xilinxmultiregimpl99_regs0;
end

always @(posedge hdmi_in1_pix2x_clk) begin
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_reset_lateness) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness <= 8'd128;
	end else begin
		if (((((~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_busy) & (~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_busy)) & (~hdmi2usbsoc_hdmi_in1_s6datacapture0_too_late)) & (~hdmi2usbsoc_hdmi_in1_s6datacapture0_too_early))) begin
			if ((hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_valid & hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_incdec)) begin
				hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness <= (hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness - 1'd1);
			end
			if ((hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_valid & (~hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_incdec))) begin
				hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness <= (hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness + 1'd1);
			end
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_pending)) begin
		if ((hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_cal | hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_ce)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_busy)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_pending)) begin
		if ((hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_cal | hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_ce)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_busy)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr <= {hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr2, hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr[9:5]};
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_i);
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_reset_lateness) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness <= 8'd128;
	end else begin
		if (((((~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_busy) & (~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_busy)) & (~hdmi2usbsoc_hdmi_in1_s6datacapture1_too_late)) & (~hdmi2usbsoc_hdmi_in1_s6datacapture1_too_early))) begin
			if ((hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_valid & hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_incdec)) begin
				hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness <= (hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness - 1'd1);
			end
			if ((hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_valid & (~hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_incdec))) begin
				hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness <= (hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness + 1'd1);
			end
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_pending)) begin
		if ((hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_cal | hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_ce)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_busy)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_pending)) begin
		if ((hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_cal | hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_ce)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_busy)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr <= {hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr2, hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr[9:5]};
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_i);
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_reset_lateness) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness <= 8'd128;
	end else begin
		if (((((~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_busy) & (~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_busy)) & (~hdmi2usbsoc_hdmi_in1_s6datacapture2_too_late)) & (~hdmi2usbsoc_hdmi_in1_s6datacapture2_too_early))) begin
			if ((hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_valid & hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_incdec)) begin
				hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness <= (hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness - 1'd1);
			end
			if ((hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_valid & (~hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_incdec))) begin
				hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness <= (hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness + 1'd1);
			end
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_pending)) begin
		if ((hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_cal | hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_ce)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_busy)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_i <= 1'd0;
	if ((~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_pending)) begin
		if ((hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_cal | hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_ce)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_pending <= 1'd1;
		end
	end else begin
		if ((~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_busy)) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_i <= 1'd1;
			hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr <= {hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr2, hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr[9:5]};
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_i);
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_o;
	if (hdmi_in1_pix2x_rst) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_lateness <= 8'd128;
		hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr <= 10'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_lateness <= 8'd128;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr <= 10'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_lateness <= 8'd128;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr <= 10'd0;
	end
	xilinxmultiregimpl56_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_i;
	xilinxmultiregimpl56_regs1 <= xilinxmultiregimpl56_regs0;
	xilinxmultiregimpl57_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_i;
	xilinxmultiregimpl57_regs1 <= xilinxmultiregimpl57_regs0;
	xilinxmultiregimpl58_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_i;
	xilinxmultiregimpl58_regs1 <= xilinxmultiregimpl58_regs0;
	xilinxmultiregimpl59_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_i;
	xilinxmultiregimpl59_regs1 <= xilinxmultiregimpl59_regs0;
	xilinxmultiregimpl60_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_i;
	xilinxmultiregimpl60_regs1 <= xilinxmultiregimpl60_regs0;
	xilinxmultiregimpl61_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_i;
	xilinxmultiregimpl61_regs1 <= xilinxmultiregimpl61_regs0;
	xilinxmultiregimpl63_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_i;
	xilinxmultiregimpl63_regs1 <= xilinxmultiregimpl63_regs0;
	xilinxmultiregimpl69_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_i;
	xilinxmultiregimpl69_regs1 <= xilinxmultiregimpl69_regs0;
	xilinxmultiregimpl70_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_i;
	xilinxmultiregimpl70_regs1 <= xilinxmultiregimpl70_regs0;
	xilinxmultiregimpl71_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_i;
	xilinxmultiregimpl71_regs1 <= xilinxmultiregimpl71_regs0;
	xilinxmultiregimpl72_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_i;
	xilinxmultiregimpl72_regs1 <= xilinxmultiregimpl72_regs0;
	xilinxmultiregimpl73_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_i;
	xilinxmultiregimpl73_regs1 <= xilinxmultiregimpl73_regs0;
	xilinxmultiregimpl74_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_i;
	xilinxmultiregimpl74_regs1 <= xilinxmultiregimpl74_regs0;
	xilinxmultiregimpl76_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_i;
	xilinxmultiregimpl76_regs1 <= xilinxmultiregimpl76_regs0;
	xilinxmultiregimpl82_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_i;
	xilinxmultiregimpl82_regs1 <= xilinxmultiregimpl82_regs0;
	xilinxmultiregimpl83_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_i;
	xilinxmultiregimpl83_regs1 <= xilinxmultiregimpl83_regs0;
	xilinxmultiregimpl84_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_i;
	xilinxmultiregimpl84_regs1 <= xilinxmultiregimpl84_regs0;
	xilinxmultiregimpl85_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_i;
	xilinxmultiregimpl85_regs1 <= xilinxmultiregimpl85_regs0;
	xilinxmultiregimpl86_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_i;
	xilinxmultiregimpl86_regs1 <= xilinxmultiregimpl86_regs0;
	xilinxmultiregimpl87_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_i;
	xilinxmultiregimpl87_regs1 <= xilinxmultiregimpl87_regs0;
	xilinxmultiregimpl89_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_i;
	xilinxmultiregimpl89_regs1 <= xilinxmultiregimpl89_regs0;
end

always @(posedge hdmi_in1_pix_o_clk) begin
	hdmi2usbsoc_hdmi_in1_syncpol_c0 <= hdmi2usbsoc_hdmi_in1_syncpol_data_in0_raw;
	hdmi2usbsoc_hdmi_in1_syncpol_c1 <= hdmi2usbsoc_hdmi_in1_syncpol_data_in1_raw;
	hdmi2usbsoc_hdmi_in1_syncpol_c2 <= hdmi2usbsoc_hdmi_in1_syncpol_data_in2_raw;
	if (hdmi_in1_pix_o_rst) begin
		hdmi2usbsoc_hdmi_in1_syncpol_c0 <= 10'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_c1 <= 10'd0;
		hdmi2usbsoc_hdmi_in1_syncpol_c2 <= 10'd0;
	end
end

always @(posedge hdmi_out0_pix_clk) begin
	hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_binary <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next_binary;
	hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q_next;
	hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_binary <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next_binary;
	hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q_next;
	if (hdmi2usbsoc_litedramportconverter0_counter_ce) begin
		hdmi2usbsoc_litedramportconverter0_counter <= (hdmi2usbsoc_litedramportconverter0_counter + 1'd1);
	end
	if ((hdmi2usbsoc_litedramportconverter0_rdata_converter_source_valid & hdmi2usbsoc_litedramportconverter0_rdata_converter_source_ready)) begin
		hdmi2usbsoc_litedramportconverter0_rdata_chunk <= {hdmi2usbsoc_litedramportconverter0_rdata_chunk[2:0], hdmi2usbsoc_litedramportconverter0_rdata_chunk[3]};
	end
	if (((hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_we & hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_writable) & (~hdmi2usbsoc_litedramportconverter0_cmd_buffer_replace))) begin
		hdmi2usbsoc_litedramportconverter0_cmd_buffer_produce <= (hdmi2usbsoc_litedramportconverter0_cmd_buffer_produce + 1'd1);
	end
	if (hdmi2usbsoc_litedramportconverter0_cmd_buffer_do_read) begin
		hdmi2usbsoc_litedramportconverter0_cmd_buffer_consume <= (hdmi2usbsoc_litedramportconverter0_cmd_buffer_consume + 1'd1);
	end
	if (((hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_we & hdmi2usbsoc_litedramportconverter0_cmd_buffer_syncfifo0_writable) & (~hdmi2usbsoc_litedramportconverter0_cmd_buffer_replace))) begin
		if ((~hdmi2usbsoc_litedramportconverter0_cmd_buffer_do_read)) begin
			hdmi2usbsoc_litedramportconverter0_cmd_buffer_level <= (hdmi2usbsoc_litedramportconverter0_cmd_buffer_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_litedramportconverter0_cmd_buffer_do_read) begin
			hdmi2usbsoc_litedramportconverter0_cmd_buffer_level <= (hdmi2usbsoc_litedramportconverter0_cmd_buffer_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_litedramportconverter0_rdata_buffer_pipe_ce) begin
		hdmi2usbsoc_litedramportconverter0_rdata_buffer_valid_n <= hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_valid;
	end
	if (hdmi2usbsoc_litedramportconverter0_rdata_buffer_pipe_ce) begin
		hdmi2usbsoc_litedramportconverter0_rdata_buffer_first_n <= (hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_valid & hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_first);
		hdmi2usbsoc_litedramportconverter0_rdata_buffer_last_n <= (hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_valid & hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_last);
	end
	if (hdmi2usbsoc_litedramportconverter0_rdata_buffer_pipe_ce) begin
		hdmi2usbsoc_litedramportconverter0_rdata_buffer_source_payload_data <= hdmi2usbsoc_litedramportconverter0_rdata_buffer_sink_payload_data;
	end
	if ((hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_valid & hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_source_ready)) begin
		if (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_last) begin
			hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_mux <= 1'd0;
		end else begin
			hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_mux <= (hdmi2usbsoc_litedramportconverter0_rdata_converter_converter_mux + 1'd1);
		end
	end
	hdmi2usbsoc_hdmi_out0_de_r <= hdmi2usbsoc_hdmi_out0_core_source_source_param_de;
	hdmi2usbsoc_hdmi_out0_core_source_valid_d <= hdmi2usbsoc_hdmi_out0_core_source_source_valid;
	hdmi2usbsoc_hdmi_out0_core_source_data_d <= hdmi2usbsoc_hdmi_out0_core_source_source_payload_data;
	if (hdmi2usbsoc_hdmi_out0_core_underflow_enable) begin
		if ((~hdmi2usbsoc_hdmi_out0_core_source_source_valid)) begin
			hdmi2usbsoc_hdmi_out0_core_underflow_counter <= (hdmi2usbsoc_hdmi_out0_core_underflow_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_out0_core_underflow_counter <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_out0_core_underflow_update) begin
		hdmi2usbsoc_hdmi_out0_core_underflow_counter_status <= hdmi2usbsoc_hdmi_out0_core_underflow_counter;
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary;
	hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q_next;
	if ((~hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_valid)) begin
		hdmi2usbsoc_hdmi_out0_core_timinggenerator_hactive <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_timinggenerator_vactive <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_ready) begin
			hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_last <= 1'd0;
			hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter <= (hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter + 1'd1);
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter == 1'd0)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_hactive <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hres)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_hactive <= 1'd0;
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hsync_start)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_hsync <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hsync_end)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_hsync <= 1'd0;
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_hscan)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_hcounter <= 1'd0;
				if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vscan)) begin
					hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter <= 1'd0;
					hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_last <= 1'd1;
				end else begin
					hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter <= (hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter + 1'd1);
				end
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter == 1'd0)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_vactive <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vres)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_vactive <= 1'd0;
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vsync_start)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_vsync <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out0_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out0_core_timinggenerator_sink_payload_vsync_end)) begin
				hdmi2usbsoc_hdmi_out0_core_timinggenerator_source_payload_vsync <= 1'd0;
			end
		end
	end
	if (hdmi2usbsoc_hdmi_out0_core_dmareader_request_issued) begin
		if ((~hdmi2usbsoc_hdmi_out0_core_dmareader_data_dequeued)) begin
			hdmi2usbsoc_hdmi_out0_core_dmareader_rsv_level <= (hdmi2usbsoc_hdmi_out0_core_dmareader_rsv_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out0_core_dmareader_data_dequeued) begin
			hdmi2usbsoc_hdmi_out0_core_dmareader_rsv_level <= (hdmi2usbsoc_hdmi_out0_core_dmareader_rsv_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_re) begin
		hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_readable <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_re) begin
			hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_readable <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_produce <= (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_consume <= (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 <= (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 <= (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_level0 - 1'd1);
		end
	end
	videoout0_state <= videoout0_next_state;
	if (hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value_ce) begin
		hdmi2usbsoc_hdmi_out0_core_dmareader_offset <= hdmi2usbsoc_hdmi_out0_core_dmareader_offset_videoout0_next_value;
	end
	hdmi2usbsoc_hdmi_out0_core_toggle_o_r <= hdmi2usbsoc_hdmi_out0_core_toggle_o;
	if ((hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out0_resetinserter_sink_sink_ready)) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_parity_in <= (~hdmi2usbsoc_hdmi_out0_resetinserter_parity_in);
	end
	if ((hdmi2usbsoc_hdmi_out0_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out0_resetinserter_source_source_ready)) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_parity_out <= (~hdmi2usbsoc_hdmi_out0_resetinserter_parity_out);
	end
	if (((hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_produce <= (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_consume <= (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level <= (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level <= (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level - 1'd1);
		end
	end
	if (((hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_produce <= (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_consume <= (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level <= (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level <= (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level - 1'd1);
		end
	end
	if (((hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_produce <= (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_consume <= (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level <= (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level <= (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_out0_resetinserter_reset) begin
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_level <= 3'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_produce <= 2'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_consume <= 2'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_level <= 3'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_produce <= 2'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_consume <= 2'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_level <= 3'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_produce <= 2'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_consume <= 2'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_parity_in <= 1'd0;
		hdmi2usbsoc_hdmi_out0_resetinserter_parity_out <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_valid_n0 <= hdmi2usbsoc_hdmi_out0_sink_valid;
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_valid_n1 <= hdmi2usbsoc_hdmi_out0_valid_n0;
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_valid_n2 <= hdmi2usbsoc_hdmi_out0_valid_n1;
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_valid_n3 <= hdmi2usbsoc_hdmi_out0_valid_n2;
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_first_n0 <= (hdmi2usbsoc_hdmi_out0_sink_valid & hdmi2usbsoc_hdmi_out0_sink_first);
		hdmi2usbsoc_hdmi_out0_last_n0 <= (hdmi2usbsoc_hdmi_out0_sink_valid & hdmi2usbsoc_hdmi_out0_sink_last);
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_first_n1 <= hdmi2usbsoc_hdmi_out0_first_n0;
		hdmi2usbsoc_hdmi_out0_last_n1 <= hdmi2usbsoc_hdmi_out0_last_n0;
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_first_n2 <= hdmi2usbsoc_hdmi_out0_first_n1;
		hdmi2usbsoc_hdmi_out0_last_n2 <= hdmi2usbsoc_hdmi_out0_last_n1;
	end
	if (hdmi2usbsoc_hdmi_out0_pipe_ce) begin
		hdmi2usbsoc_hdmi_out0_first_n3 <= hdmi2usbsoc_hdmi_out0_first_n2;
		hdmi2usbsoc_hdmi_out0_last_n3 <= hdmi2usbsoc_hdmi_out0_last_n2;
	end
	if (hdmi2usbsoc_hdmi_out0_ce) begin
		hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_y <= hdmi2usbsoc_hdmi_out0_sink_y;
		hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out0_sink_cb;
		hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out0_sink_cr;
		hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_y <= hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_y;
		hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_y <= hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_y;
		hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out0_record1_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_out0_record3_ycbcr_n_y <= hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_y;
		hdmi2usbsoc_hdmi_out0_record3_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_out0_record3_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out0_record2_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_out0_cb_minus_coffset <= (hdmi2usbsoc_hdmi_out0_sink_cb - 8'd128);
		hdmi2usbsoc_hdmi_out0_cr_minus_coffset <= (hdmi2usbsoc_hdmi_out0_sink_cr - 8'd128);
		hdmi2usbsoc_hdmi_out0_y_minus_yoffset <= (hdmi2usbsoc_hdmi_out0_record0_ycbcr_n_y - 5'd16);
		hdmi2usbsoc_hdmi_out0_cr_minus_coffset_mult_acoef <= (hdmi2usbsoc_hdmi_out0_cr_minus_coffset * $signed({1'd0, 7'd98}));
		hdmi2usbsoc_hdmi_out0_cb_minus_coffset_mult_bcoef <= (hdmi2usbsoc_hdmi_out0_cb_minus_coffset * 5'sd23);
		hdmi2usbsoc_hdmi_out0_cr_minus_coffset_mult_ccoef <= (hdmi2usbsoc_hdmi_out0_cr_minus_coffset * 6'sd41);
		hdmi2usbsoc_hdmi_out0_cb_minus_coffset_mult_dcoef <= (hdmi2usbsoc_hdmi_out0_cb_minus_coffset * $signed({1'd0, 7'd116}));
		hdmi2usbsoc_hdmi_out0_r <= (hdmi2usbsoc_hdmi_out0_y_minus_yoffset + hdmi2usbsoc_hdmi_out0_cr_minus_coffset_mult_acoef[19:6]);
		hdmi2usbsoc_hdmi_out0_g <= ((hdmi2usbsoc_hdmi_out0_y_minus_yoffset + hdmi2usbsoc_hdmi_out0_cb_minus_coffset_mult_bcoef[19:6]) + hdmi2usbsoc_hdmi_out0_cr_minus_coffset_mult_ccoef[19:6]);
		hdmi2usbsoc_hdmi_out0_b <= (hdmi2usbsoc_hdmi_out0_y_minus_yoffset + hdmi2usbsoc_hdmi_out0_cb_minus_coffset_mult_dcoef[19:6]);
		if ((hdmi2usbsoc_hdmi_out0_r > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_out0_source_r <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_out0_r < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_out0_source_r <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_out0_source_r <= hdmi2usbsoc_hdmi_out0_r;
			end
		end
		if ((hdmi2usbsoc_hdmi_out0_g > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_out0_source_g <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_out0_g < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_out0_source_g <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_out0_source_g <= hdmi2usbsoc_hdmi_out0_g;
			end
		end
		if ((hdmi2usbsoc_hdmi_out0_b > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_out0_source_b <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_out0_b < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_out0_source_b <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_out0_source_b <= hdmi2usbsoc_hdmi_out0_b;
			end
		end
	end
	hdmi2usbsoc_hdmi_out0_next_s0 <= hdmi2usbsoc_hdmi_out0_sink_payload_hsync;
	hdmi2usbsoc_hdmi_out0_next_s1 <= hdmi2usbsoc_hdmi_out0_next_s0;
	hdmi2usbsoc_hdmi_out0_next_s2 <= hdmi2usbsoc_hdmi_out0_next_s1;
	hdmi2usbsoc_hdmi_out0_next_s3 <= hdmi2usbsoc_hdmi_out0_next_s2;
	hdmi2usbsoc_hdmi_out0_next_s4 <= hdmi2usbsoc_hdmi_out0_next_s3;
	hdmi2usbsoc_hdmi_out0_next_s5 <= hdmi2usbsoc_hdmi_out0_next_s4;
	hdmi2usbsoc_hdmi_out0_next_s6 <= hdmi2usbsoc_hdmi_out0_sink_payload_vsync;
	hdmi2usbsoc_hdmi_out0_next_s7 <= hdmi2usbsoc_hdmi_out0_next_s6;
	hdmi2usbsoc_hdmi_out0_next_s8 <= hdmi2usbsoc_hdmi_out0_next_s7;
	hdmi2usbsoc_hdmi_out0_next_s9 <= hdmi2usbsoc_hdmi_out0_next_s8;
	hdmi2usbsoc_hdmi_out0_next_s10 <= hdmi2usbsoc_hdmi_out0_next_s9;
	hdmi2usbsoc_hdmi_out0_next_s11 <= hdmi2usbsoc_hdmi_out0_next_s10;
	hdmi2usbsoc_hdmi_out0_next_s12 <= hdmi2usbsoc_hdmi_out0_sink_payload_de;
	hdmi2usbsoc_hdmi_out0_next_s13 <= hdmi2usbsoc_hdmi_out0_next_s12;
	hdmi2usbsoc_hdmi_out0_next_s14 <= hdmi2usbsoc_hdmi_out0_next_s13;
	hdmi2usbsoc_hdmi_out0_next_s15 <= hdmi2usbsoc_hdmi_out0_next_s14;
	hdmi2usbsoc_hdmi_out0_next_s16 <= hdmi2usbsoc_hdmi_out0_next_s15;
	hdmi2usbsoc_hdmi_out0_next_s17 <= hdmi2usbsoc_hdmi_out0_next_s16;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1d <= (((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[0] + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[1]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[2]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[3]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[4]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[5]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[6]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0[7]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0];
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[1] <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[2] <= ((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[3] <= ((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[4] <= ((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[5] <= ((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[6] <= ((((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[6]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[7] <= ((((((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[6]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_d1[7]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[8] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m <= ((((((((~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[0]) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[1])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[2])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[3])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[4])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[5])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[6])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[7]));
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m <= (((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[0] + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[1]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[2]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[3]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[4]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[5]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[6]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m[7]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c0 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_c;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de0 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_de;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c2 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_c1;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de2 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de1;
	if (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_new_de2) begin
		if (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m == hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m)}))) begin
			hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[9] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]);
			hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
			if (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]) begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m}));
			end
		end else begin
			if ((((~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt[5]) & $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m > hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m)})) | (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt[5] & $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m > hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m)})))) begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[9] <= 1'd1;
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt <= (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, {hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[9] <= 1'd0;
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt <= (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt - $signed({1'd0, {(~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_n0q_m}));
			end
		end
	end else begin
		hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out <= sync_f_array_muxed0;
		hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cnt <= 1'd0;
	end
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1d <= (((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[0] + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[1]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[2]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[3]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[4]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[5]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[6]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0[7]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0];
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[1] <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[2] <= ((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[3] <= ((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[4] <= ((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[5] <= ((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[6] <= ((((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[6]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[7] <= ((((((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[6]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_d1[7]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[8] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m <= ((((((((~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[0]) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[1])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[2])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[3])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[4])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[5])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[6])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[7]));
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m <= (((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[0] + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[1]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[2]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[3]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[4]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[5]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[6]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m[7]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c0 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_c;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de0 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_de;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c2 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_c1;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de2 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de1;
	if (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_new_de2) begin
		if (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m == hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m)}))) begin
			hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[9] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]);
			hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
			if (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]) begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m}));
			end
		end else begin
			if ((((~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt[5]) & $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m > hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m)})) | (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt[5] & $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m > hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m)})))) begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[9] <= 1'd1;
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt <= (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, {hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[9] <= 1'd0;
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt <= (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt - $signed({1'd0, {(~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_n0q_m}));
			end
		end
	end else begin
		hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out <= sync_f_array_muxed1;
		hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cnt <= 1'd0;
	end
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1d <= (((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[0] + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[1]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[2]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[3]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[4]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[5]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[6]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0[7]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0];
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[1] <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[2] <= ((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[3] <= ((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[4] <= ((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[5] <= ((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[6] <= ((((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[6]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[7] <= ((((((((((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[6]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_d1[7]) ^ hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[8] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m <= ((((((((~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[0]) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[1])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[2])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[3])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[4])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[5])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[6])) + (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[7]));
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m <= (((((((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[0] + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[1]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[2]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[3]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[4]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[5]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[6]) + hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m[7]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c0 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_c;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de0 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_de;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de1 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de0;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c2 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_c1;
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de2 <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de1;
	if (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_new_de2) begin
		if (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m == hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m)}))) begin
			hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[9] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]);
			hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
			if (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]) begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt <= ((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m}));
			end
		end else begin
			if ((((~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt[5]) & $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m > hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m)})) | (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt[5] & $signed({1'd0, (hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m > hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m)})))) begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[9] <= 1'd1;
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= (~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt <= (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, {hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[9] <= 1'd0;
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[8] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt <= (((hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt - $signed({1'd0, {(~hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_n0q_m}));
			end
		end
	end else begin
		hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out <= sync_f_array_muxed2;
		hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cnt <= 1'd0;
	end
	xilinxmultiregimpl102_regs0 <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q;
	xilinxmultiregimpl102_regs1 <= xilinxmultiregimpl102_regs0;
	xilinxmultiregimpl103_regs0 <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q;
	xilinxmultiregimpl103_regs1 <= xilinxmultiregimpl103_regs0;
	xilinxmultiregimpl105_regs0 <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q;
	xilinxmultiregimpl105_regs1 <= xilinxmultiregimpl105_regs0;
	xilinxmultiregimpl108_regs0 <= hdmi2usbsoc_hdmi_out0_core_toggle_i;
	xilinxmultiregimpl108_regs1 <= xilinxmultiregimpl108_regs0;
end

always @(posedge hdmi_out0_pix2x_clk) begin
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x_pol <= (hdmi_out0_pix_clk ? hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[4:0] : hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_out[9:5]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x_pol <= (hdmi_out0_pix_clk ? hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[4:0] : hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_out[9:5]);
	hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x_pol <= (hdmi_out0_pix_clk ? hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[4:0] : hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_out[9:5]);
end

always @(posedge hdmi_out1_pix_clk) begin
	hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_binary <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next_binary;
	hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q_next;
	hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_binary <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next_binary;
	hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q_next;
	if (hdmi2usbsoc_litedramportconverter1_counter_ce) begin
		hdmi2usbsoc_litedramportconverter1_counter <= (hdmi2usbsoc_litedramportconverter1_counter + 1'd1);
	end
	if ((hdmi2usbsoc_litedramportconverter1_rdata_converter_source_valid & hdmi2usbsoc_litedramportconverter1_rdata_converter_source_ready)) begin
		hdmi2usbsoc_litedramportconverter1_rdata_chunk <= {hdmi2usbsoc_litedramportconverter1_rdata_chunk[2:0], hdmi2usbsoc_litedramportconverter1_rdata_chunk[3]};
	end
	if (((hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_we & hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_writable) & (~hdmi2usbsoc_litedramportconverter1_cmd_buffer_replace))) begin
		hdmi2usbsoc_litedramportconverter1_cmd_buffer_produce <= (hdmi2usbsoc_litedramportconverter1_cmd_buffer_produce + 1'd1);
	end
	if (hdmi2usbsoc_litedramportconverter1_cmd_buffer_do_read) begin
		hdmi2usbsoc_litedramportconverter1_cmd_buffer_consume <= (hdmi2usbsoc_litedramportconverter1_cmd_buffer_consume + 1'd1);
	end
	if (((hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_we & hdmi2usbsoc_litedramportconverter1_cmd_buffer_syncfifo1_writable) & (~hdmi2usbsoc_litedramportconverter1_cmd_buffer_replace))) begin
		if ((~hdmi2usbsoc_litedramportconverter1_cmd_buffer_do_read)) begin
			hdmi2usbsoc_litedramportconverter1_cmd_buffer_level <= (hdmi2usbsoc_litedramportconverter1_cmd_buffer_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_litedramportconverter1_cmd_buffer_do_read) begin
			hdmi2usbsoc_litedramportconverter1_cmd_buffer_level <= (hdmi2usbsoc_litedramportconverter1_cmd_buffer_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_litedramportconverter1_rdata_buffer_pipe_ce) begin
		hdmi2usbsoc_litedramportconverter1_rdata_buffer_valid_n <= hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_valid;
	end
	if (hdmi2usbsoc_litedramportconverter1_rdata_buffer_pipe_ce) begin
		hdmi2usbsoc_litedramportconverter1_rdata_buffer_first_n <= (hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_valid & hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_first);
		hdmi2usbsoc_litedramportconverter1_rdata_buffer_last_n <= (hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_valid & hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_last);
	end
	if (hdmi2usbsoc_litedramportconverter1_rdata_buffer_pipe_ce) begin
		hdmi2usbsoc_litedramportconverter1_rdata_buffer_source_payload_data <= hdmi2usbsoc_litedramportconverter1_rdata_buffer_sink_payload_data;
	end
	if ((hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_valid & hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_source_ready)) begin
		if (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_last) begin
			hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_mux <= 1'd0;
		end else begin
			hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_mux <= (hdmi2usbsoc_litedramportconverter1_rdata_converter_converter_mux + 1'd1);
		end
	end
	hdmi2usbsoc_hdmi_out1_de_r <= hdmi2usbsoc_hdmi_out1_core_source_source_param_de;
	hdmi2usbsoc_hdmi_out1_core_source_valid_d <= hdmi2usbsoc_hdmi_out1_core_source_source_valid;
	hdmi2usbsoc_hdmi_out1_core_source_data_d <= hdmi2usbsoc_hdmi_out1_core_source_source_payload_data;
	if (hdmi2usbsoc_hdmi_out1_core_underflow_enable) begin
		if ((~hdmi2usbsoc_hdmi_out1_core_source_source_valid)) begin
			hdmi2usbsoc_hdmi_out1_core_underflow_counter <= (hdmi2usbsoc_hdmi_out1_core_underflow_counter + 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi_out1_core_underflow_counter <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_out1_core_underflow_update) begin
		hdmi2usbsoc_hdmi_out1_core_underflow_counter_status <= hdmi2usbsoc_hdmi_out1_core_underflow_counter;
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_binary <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next_binary;
	hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q_next;
	if ((~hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_valid)) begin
		hdmi2usbsoc_hdmi_out1_core_timinggenerator_hactive <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_timinggenerator_vactive <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_ready) begin
			hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_last <= 1'd0;
			hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter <= (hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter + 1'd1);
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter == 1'd0)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_hactive <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hres)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_hactive <= 1'd0;
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hsync_start)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_hsync <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hsync_end)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_hsync <= 1'd0;
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_hscan)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_hcounter <= 1'd0;
				if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vscan)) begin
					hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter <= 1'd0;
					hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_last <= 1'd1;
				end else begin
					hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter <= (hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter + 1'd1);
				end
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter == 1'd0)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_vactive <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vres)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_vactive <= 1'd0;
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vsync_start)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_vsync <= 1'd1;
			end
			if ((hdmi2usbsoc_hdmi_out1_core_timinggenerator_vcounter == hdmi2usbsoc_hdmi_out1_core_timinggenerator_sink_payload_vsync_end)) begin
				hdmi2usbsoc_hdmi_out1_core_timinggenerator_source_payload_vsync <= 1'd0;
			end
		end
	end
	if (hdmi2usbsoc_hdmi_out1_core_dmareader_request_issued) begin
		if ((~hdmi2usbsoc_hdmi_out1_core_dmareader_data_dequeued)) begin
			hdmi2usbsoc_hdmi_out1_core_dmareader_rsv_level <= (hdmi2usbsoc_hdmi_out1_core_dmareader_rsv_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out1_core_dmareader_data_dequeued) begin
			hdmi2usbsoc_hdmi_out1_core_dmareader_rsv_level <= (hdmi2usbsoc_hdmi_out1_core_dmareader_rsv_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_re) begin
		hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_readable <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_re) begin
			hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_readable <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_produce <= (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_consume <= (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 <= (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 <= (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_level0 - 1'd1);
		end
	end
	videoout1_state <= videoout1_next_state;
	if (hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value_ce) begin
		hdmi2usbsoc_hdmi_out1_core_dmareader_offset <= hdmi2usbsoc_hdmi_out1_core_dmareader_offset_videoout1_next_value;
	end
	hdmi2usbsoc_hdmi_out1_core_toggle_o_r <= hdmi2usbsoc_hdmi_out1_core_toggle_o;
	if ((hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_valid & hdmi2usbsoc_hdmi_out1_resetinserter_sink_sink_ready)) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_parity_in <= (~hdmi2usbsoc_hdmi_out1_resetinserter_parity_in);
	end
	if ((hdmi2usbsoc_hdmi_out1_resetinserter_source_source_valid & hdmi2usbsoc_hdmi_out1_resetinserter_source_source_ready)) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_parity_out <= (~hdmi2usbsoc_hdmi_out1_resetinserter_parity_out);
	end
	if (((hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_produce <= (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_consume <= (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level <= (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level <= (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level - 1'd1);
		end
	end
	if (((hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_produce <= (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_consume <= (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level <= (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level <= (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level - 1'd1);
		end
	end
	if (((hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_replace))) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_produce <= (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_do_read) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_consume <= (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_we & hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level <= (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_do_read) begin
			hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level <= (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_out1_resetinserter_reset) begin
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_level <= 3'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_produce <= 2'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_consume <= 2'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_level <= 3'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_produce <= 2'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_consume <= 2'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_level <= 3'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_produce <= 2'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_consume <= 2'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_parity_in <= 1'd0;
		hdmi2usbsoc_hdmi_out1_resetinserter_parity_out <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_valid_n0 <= hdmi2usbsoc_hdmi_out1_sink_valid;
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_valid_n1 <= hdmi2usbsoc_hdmi_out1_valid_n0;
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_valid_n2 <= hdmi2usbsoc_hdmi_out1_valid_n1;
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_valid_n3 <= hdmi2usbsoc_hdmi_out1_valid_n2;
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_first_n0 <= (hdmi2usbsoc_hdmi_out1_sink_valid & hdmi2usbsoc_hdmi_out1_sink_first);
		hdmi2usbsoc_hdmi_out1_last_n0 <= (hdmi2usbsoc_hdmi_out1_sink_valid & hdmi2usbsoc_hdmi_out1_sink_last);
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_first_n1 <= hdmi2usbsoc_hdmi_out1_first_n0;
		hdmi2usbsoc_hdmi_out1_last_n1 <= hdmi2usbsoc_hdmi_out1_last_n0;
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_first_n2 <= hdmi2usbsoc_hdmi_out1_first_n1;
		hdmi2usbsoc_hdmi_out1_last_n2 <= hdmi2usbsoc_hdmi_out1_last_n1;
	end
	if (hdmi2usbsoc_hdmi_out1_pipe_ce) begin
		hdmi2usbsoc_hdmi_out1_first_n3 <= hdmi2usbsoc_hdmi_out1_first_n2;
		hdmi2usbsoc_hdmi_out1_last_n3 <= hdmi2usbsoc_hdmi_out1_last_n2;
	end
	if (hdmi2usbsoc_hdmi_out1_ce) begin
		hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_y <= hdmi2usbsoc_hdmi_out1_sink_y;
		hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out1_sink_cb;
		hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out1_sink_cr;
		hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_y <= hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_y;
		hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_y <= hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_y;
		hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out1_record1_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_out1_record3_ycbcr_n_y <= hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_y;
		hdmi2usbsoc_hdmi_out1_record3_ycbcr_n_cb <= hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_cb;
		hdmi2usbsoc_hdmi_out1_record3_ycbcr_n_cr <= hdmi2usbsoc_hdmi_out1_record2_ycbcr_n_cr;
		hdmi2usbsoc_hdmi_out1_cb_minus_coffset <= (hdmi2usbsoc_hdmi_out1_sink_cb - 8'd128);
		hdmi2usbsoc_hdmi_out1_cr_minus_coffset <= (hdmi2usbsoc_hdmi_out1_sink_cr - 8'd128);
		hdmi2usbsoc_hdmi_out1_y_minus_yoffset <= (hdmi2usbsoc_hdmi_out1_record0_ycbcr_n_y - 5'd16);
		hdmi2usbsoc_hdmi_out1_cr_minus_coffset_mult_acoef <= (hdmi2usbsoc_hdmi_out1_cr_minus_coffset * $signed({1'd0, 7'd98}));
		hdmi2usbsoc_hdmi_out1_cb_minus_coffset_mult_bcoef <= (hdmi2usbsoc_hdmi_out1_cb_minus_coffset * 5'sd23);
		hdmi2usbsoc_hdmi_out1_cr_minus_coffset_mult_ccoef <= (hdmi2usbsoc_hdmi_out1_cr_minus_coffset * 6'sd41);
		hdmi2usbsoc_hdmi_out1_cb_minus_coffset_mult_dcoef <= (hdmi2usbsoc_hdmi_out1_cb_minus_coffset * $signed({1'd0, 7'd116}));
		hdmi2usbsoc_hdmi_out1_r <= (hdmi2usbsoc_hdmi_out1_y_minus_yoffset + hdmi2usbsoc_hdmi_out1_cr_minus_coffset_mult_acoef[19:6]);
		hdmi2usbsoc_hdmi_out1_g <= ((hdmi2usbsoc_hdmi_out1_y_minus_yoffset + hdmi2usbsoc_hdmi_out1_cb_minus_coffset_mult_bcoef[19:6]) + hdmi2usbsoc_hdmi_out1_cr_minus_coffset_mult_ccoef[19:6]);
		hdmi2usbsoc_hdmi_out1_b <= (hdmi2usbsoc_hdmi_out1_y_minus_yoffset + hdmi2usbsoc_hdmi_out1_cb_minus_coffset_mult_dcoef[19:6]);
		if ((hdmi2usbsoc_hdmi_out1_r > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_out1_source_r <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_out1_r < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_out1_source_r <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_out1_source_r <= hdmi2usbsoc_hdmi_out1_r;
			end
		end
		if ((hdmi2usbsoc_hdmi_out1_g > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_out1_source_g <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_out1_g < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_out1_source_g <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_out1_source_g <= hdmi2usbsoc_hdmi_out1_g;
			end
		end
		if ((hdmi2usbsoc_hdmi_out1_b > $signed({1'd0, 8'd255}))) begin
			hdmi2usbsoc_hdmi_out1_source_b <= 8'd255;
		end else begin
			if ((hdmi2usbsoc_hdmi_out1_b < $signed({1'd0, 1'd0}))) begin
				hdmi2usbsoc_hdmi_out1_source_b <= 1'd0;
			end else begin
				hdmi2usbsoc_hdmi_out1_source_b <= hdmi2usbsoc_hdmi_out1_b;
			end
		end
	end
	hdmi2usbsoc_hdmi_out1_next_s0 <= hdmi2usbsoc_hdmi_out1_sink_payload_hsync;
	hdmi2usbsoc_hdmi_out1_next_s1 <= hdmi2usbsoc_hdmi_out1_next_s0;
	hdmi2usbsoc_hdmi_out1_next_s2 <= hdmi2usbsoc_hdmi_out1_next_s1;
	hdmi2usbsoc_hdmi_out1_next_s3 <= hdmi2usbsoc_hdmi_out1_next_s2;
	hdmi2usbsoc_hdmi_out1_next_s4 <= hdmi2usbsoc_hdmi_out1_next_s3;
	hdmi2usbsoc_hdmi_out1_next_s5 <= hdmi2usbsoc_hdmi_out1_next_s4;
	hdmi2usbsoc_hdmi_out1_next_s6 <= hdmi2usbsoc_hdmi_out1_sink_payload_vsync;
	hdmi2usbsoc_hdmi_out1_next_s7 <= hdmi2usbsoc_hdmi_out1_next_s6;
	hdmi2usbsoc_hdmi_out1_next_s8 <= hdmi2usbsoc_hdmi_out1_next_s7;
	hdmi2usbsoc_hdmi_out1_next_s9 <= hdmi2usbsoc_hdmi_out1_next_s8;
	hdmi2usbsoc_hdmi_out1_next_s10 <= hdmi2usbsoc_hdmi_out1_next_s9;
	hdmi2usbsoc_hdmi_out1_next_s11 <= hdmi2usbsoc_hdmi_out1_next_s10;
	hdmi2usbsoc_hdmi_out1_next_s12 <= hdmi2usbsoc_hdmi_out1_sink_payload_de;
	hdmi2usbsoc_hdmi_out1_next_s13 <= hdmi2usbsoc_hdmi_out1_next_s12;
	hdmi2usbsoc_hdmi_out1_next_s14 <= hdmi2usbsoc_hdmi_out1_next_s13;
	hdmi2usbsoc_hdmi_out1_next_s15 <= hdmi2usbsoc_hdmi_out1_next_s14;
	hdmi2usbsoc_hdmi_out1_next_s16 <= hdmi2usbsoc_hdmi_out1_next_s15;
	hdmi2usbsoc_hdmi_out1_next_s17 <= hdmi2usbsoc_hdmi_out1_next_s16;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1d <= (((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[0] + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[1]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[2]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[3]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[4]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[5]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[6]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0[7]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0];
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[1] <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[2] <= ((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[3] <= ((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[4] <= ((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[5] <= ((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[6] <= ((((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[6]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[7] <= ((((((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[6]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_d1[7]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[8] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m <= ((((((((~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[0]) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[1])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[2])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[3])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[4])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[5])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[6])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[7]));
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m <= (((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[0] + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[1]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[2]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[3]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[4]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[5]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[6]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m[7]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c0 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_c;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de0 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_de;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c2 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_c1;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de2 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de1;
	if (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_new_de2) begin
		if (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m == hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m)}))) begin
			hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[9] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[8]);
			hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[8];
			if (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[8]) begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[7:0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[7:0] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m}));
			end
		end else begin
			if ((((~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt[5]) & $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m > hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m)})) | (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt[5] & $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m > hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m)})))) begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[9] <= 1'd1;
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[8];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[7:0] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt <= (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt + $signed({1'd0, {hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[9] <= 1'd0;
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[8];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[7:0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt <= (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt - $signed({1'd0, {(~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_n0q_m}));
			end
		end
	end else begin
		hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out <= sync_f_array_muxed3;
		hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cnt <= 1'd0;
	end
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1d <= (((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[0] + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[1]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[2]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[3]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[4]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[5]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[6]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0[7]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0];
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[1] <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[2] <= ((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[3] <= ((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[4] <= ((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[5] <= ((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[6] <= ((((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[6]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[7] <= ((((((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[6]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_d1[7]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[8] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m <= ((((((((~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[0]) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[1])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[2])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[3])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[4])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[5])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[6])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[7]));
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m <= (((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[0] + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[1]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[2]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[3]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[4]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[5]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[6]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m[7]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c0 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_c;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de0 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_de;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c2 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_c1;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de2 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de1;
	if (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_new_de2) begin
		if (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m == hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m)}))) begin
			hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[9] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[8]);
			hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[8];
			if (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[8]) begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[7:0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[7:0] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m}));
			end
		end else begin
			if ((((~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt[5]) & $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m > hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m)})) | (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt[5] & $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m > hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m)})))) begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[9] <= 1'd1;
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[8];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[7:0] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt <= (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt + $signed({1'd0, {hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[9] <= 1'd0;
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[8];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[7:0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt <= (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt - $signed({1'd0, {(~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_n0q_m}));
			end
		end
	end else begin
		hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out <= sync_f_array_muxed4;
		hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cnt <= 1'd0;
	end
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1d <= (((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[0] + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[1]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[2]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[3]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[4]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[5]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[6]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0[7]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0];
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[1] <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[2] <= ((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[3] <= ((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[4] <= ((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[5] <= ((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[6] <= ((((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[6]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[7] <= ((((((((((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[0] ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[1]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[2]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[3]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[4]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[5]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[6]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_d1[7]) ^ hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[8] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m8_n);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m <= ((((((((~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[0]) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[1])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[2])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[3])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[4])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[5])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[6])) + (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[7]));
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m <= (((((((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[0] + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[1]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[2]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[3]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[4]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[5]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[6]) + hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m[7]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c0 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_c;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de0 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_de;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de1 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de0;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c2 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_c1;
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de2 <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de1;
	if (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_new_de2) begin
		if (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m == hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m)}))) begin
			hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[9] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[8]);
			hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[8];
			if (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[8]) begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[7:0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[7:0] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt <= ((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m}));
			end
		end else begin
			if ((((~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt[5]) & $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m > hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m)})) | (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt[5] & $signed({1'd0, (hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m > hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m)})))) begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[9] <= 1'd1;
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[8];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[7:0] <= (~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[7:0]);
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt <= (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt + $signed({1'd0, {hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[8], 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m}));
			end else begin
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[9] <= 1'd0;
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[8] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[8];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[7:0] <= hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[7:0];
				hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt <= (((hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt - $signed({1'd0, {(~hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_q_m_r[8]), 1'd0}})) + $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_n0q_m}));
			end
		end
	end else begin
		hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out <= sync_f_array_muxed5;
		hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cnt <= 1'd0;
	end
	xilinxmultiregimpl111_regs0 <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q;
	xilinxmultiregimpl111_regs1 <= xilinxmultiregimpl111_regs0;
	xilinxmultiregimpl112_regs0 <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q;
	xilinxmultiregimpl112_regs1 <= xilinxmultiregimpl112_regs0;
	xilinxmultiregimpl114_regs0 <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q;
	xilinxmultiregimpl114_regs1 <= xilinxmultiregimpl114_regs0;
	xilinxmultiregimpl117_regs0 <= hdmi2usbsoc_hdmi_out1_core_toggle_i;
	xilinxmultiregimpl117_regs1 <= xilinxmultiregimpl117_regs0;
end

always @(posedge hdmi_out1_pix2x_clk) begin
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x_pol <= (hdmi_out1_pix_clk ? hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[4:0] : hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_out[9:5]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x_pol <= (hdmi_out1_pix_clk ? hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[4:0] : hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_out[9:5]);
	hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x_pol <= (hdmi_out1_pix_clk ? hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[4:0] : hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_out[9:5]);
end

always @(posedge por_clk) begin
	if ((hdmi2usbsoc_crg_por != 1'd0)) begin
		hdmi2usbsoc_crg_por <= (hdmi2usbsoc_crg_por - 1'd1);
	end
	if (por_rst) begin
		hdmi2usbsoc_crg_por <= 11'd2047;
	end
end

always @(posedge sdram_half_clk) begin
	if ((hdmi2usbsoc_ddrphy_phase_half == hdmi2usbsoc_ddrphy_phase_sys)) begin
		hdmi2usbsoc_ddrphy_phase_sel <= 1'd0;
	end else begin
		hdmi2usbsoc_ddrphy_phase_sel <= (hdmi2usbsoc_ddrphy_phase_sel + 1'd1);
	end
	hdmi2usbsoc_ddrphy_phase_half <= (hdmi2usbsoc_ddrphy_phase_half + 1'd1);
	hdmi2usbsoc_ddrphy_record0_reset_n <= hdmi2usbsoc_ddrphy_dfi_p0_reset_n;
	hdmi2usbsoc_ddrphy_record0_odt <= hdmi2usbsoc_ddrphy_dfi_p0_odt;
	hdmi2usbsoc_ddrphy_record0_address <= hdmi2usbsoc_ddrphy_dfi_p0_address;
	hdmi2usbsoc_ddrphy_record0_bank <= hdmi2usbsoc_ddrphy_dfi_p0_bank;
	hdmi2usbsoc_ddrphy_record0_cs_n <= hdmi2usbsoc_ddrphy_dfi_p0_cs_n;
	hdmi2usbsoc_ddrphy_record0_cke <= hdmi2usbsoc_ddrphy_dfi_p0_cke;
	hdmi2usbsoc_ddrphy_record0_cas_n <= hdmi2usbsoc_ddrphy_dfi_p0_cas_n;
	hdmi2usbsoc_ddrphy_record0_ras_n <= hdmi2usbsoc_ddrphy_dfi_p0_ras_n;
	hdmi2usbsoc_ddrphy_record0_we_n <= hdmi2usbsoc_ddrphy_dfi_p0_we_n;
	hdmi2usbsoc_ddrphy_record1_reset_n <= hdmi2usbsoc_ddrphy_dfi_p1_reset_n;
	hdmi2usbsoc_ddrphy_record1_odt <= hdmi2usbsoc_ddrphy_dfi_p1_odt;
	hdmi2usbsoc_ddrphy_record1_address <= hdmi2usbsoc_ddrphy_dfi_p1_address;
	hdmi2usbsoc_ddrphy_record1_bank <= hdmi2usbsoc_ddrphy_dfi_p1_bank;
	hdmi2usbsoc_ddrphy_record1_cs_n <= hdmi2usbsoc_ddrphy_dfi_p1_cs_n;
	hdmi2usbsoc_ddrphy_record1_cke <= hdmi2usbsoc_ddrphy_dfi_p1_cke;
	hdmi2usbsoc_ddrphy_record1_cas_n <= hdmi2usbsoc_ddrphy_dfi_p1_cas_n;
	hdmi2usbsoc_ddrphy_record1_ras_n <= hdmi2usbsoc_ddrphy_dfi_p1_ras_n;
	hdmi2usbsoc_ddrphy_record1_we_n <= hdmi2usbsoc_ddrphy_dfi_p1_we_n;
	ddram_a <= sync_rhs_array_muxed0;
	ddram_ba <= sync_rhs_array_muxed1;
	ddram_cke <= sync_rhs_array_muxed2;
	ddram_ras_n <= sync_rhs_array_muxed3;
	ddram_cas_n <= sync_rhs_array_muxed4;
	ddram_we_n <= sync_rhs_array_muxed5;
	ddram_odt <= sync_rhs_array_muxed6;
	hdmi2usbsoc_ddrphy_postamble <= hdmi2usbsoc_ddrphy_drive_dqs;
	hdmi2usbsoc_ddrphy_r_dfi_wrdata_en <= {hdmi2usbsoc_ddrphy_r_dfi_wrdata_en, hdmi2usbsoc_ddrphy_wrdata_en_d};
	if (sdram_half_rst) begin
		ddram_cke <= 1'd0;
		ddram_ras_n <= 1'd0;
		ddram_cas_n <= 1'd0;
		ddram_we_n <= 1'd0;
		ddram_ba <= 3'd0;
		ddram_a <= 13'd0;
		ddram_odt <= 1'd0;
		hdmi2usbsoc_ddrphy_phase_sel <= 1'd0;
		hdmi2usbsoc_ddrphy_phase_half <= 1'd0;
		hdmi2usbsoc_ddrphy_record0_address <= 13'd0;
		hdmi2usbsoc_ddrphy_record0_bank <= 3'd0;
		hdmi2usbsoc_ddrphy_record0_cas_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record0_cs_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record0_ras_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record0_we_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record0_cke <= 1'd0;
		hdmi2usbsoc_ddrphy_record0_odt <= 1'd0;
		hdmi2usbsoc_ddrphy_record0_reset_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record1_address <= 13'd0;
		hdmi2usbsoc_ddrphy_record1_bank <= 3'd0;
		hdmi2usbsoc_ddrphy_record1_cas_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record1_cs_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record1_ras_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record1_we_n <= 1'd0;
		hdmi2usbsoc_ddrphy_record1_cke <= 1'd0;
		hdmi2usbsoc_ddrphy_record1_odt <= 1'd0;
		hdmi2usbsoc_ddrphy_record1_reset_n <= 1'd0;
		hdmi2usbsoc_ddrphy_postamble <= 1'd0;
		hdmi2usbsoc_ddrphy_r_dfi_wrdata_en <= 3'd0;
	end
end

always @(posedge sys_clk) begin
	hdmi2usbsoc_hdmi2usbsoc_rom_bus_ack <= 1'd0;
	if (((hdmi2usbsoc_hdmi2usbsoc_rom_bus_cyc & hdmi2usbsoc_hdmi2usbsoc_rom_bus_stb) & (~hdmi2usbsoc_hdmi2usbsoc_rom_bus_ack))) begin
		hdmi2usbsoc_hdmi2usbsoc_rom_bus_ack <= 1'd1;
	end
	hdmi2usbsoc_hdmi2usbsoc_sram_bus_ack <= 1'd0;
	if (((hdmi2usbsoc_hdmi2usbsoc_sram_bus_cyc & hdmi2usbsoc_hdmi2usbsoc_sram_bus_stb) & (~hdmi2usbsoc_hdmi2usbsoc_sram_bus_ack))) begin
		hdmi2usbsoc_hdmi2usbsoc_sram_bus_ack <= 1'd1;
	end
	hdmi2usbsoc_hdmi2usbsoc_interface_we <= 1'd0;
	hdmi2usbsoc_hdmi2usbsoc_interface_dat_w <= hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_dat_w;
	hdmi2usbsoc_hdmi2usbsoc_interface_adr <= hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_adr;
	hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_dat_r <= hdmi2usbsoc_hdmi2usbsoc_interface_dat_r;
	if ((hdmi2usbsoc_hdmi2usbsoc_counter == 1'd1)) begin
		hdmi2usbsoc_hdmi2usbsoc_interface_we <= hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_we;
	end
	if ((hdmi2usbsoc_hdmi2usbsoc_counter == 2'd2)) begin
		hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_ack <= 1'd1;
	end
	if ((hdmi2usbsoc_hdmi2usbsoc_counter == 2'd3)) begin
		hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_ack <= 1'd0;
	end
	if ((hdmi2usbsoc_hdmi2usbsoc_counter != 1'd0)) begin
		hdmi2usbsoc_hdmi2usbsoc_counter <= (hdmi2usbsoc_hdmi2usbsoc_counter + 1'd1);
	end else begin
		if ((hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_cyc & hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_stb)) begin
			hdmi2usbsoc_hdmi2usbsoc_counter <= 1'd1;
		end
	end
	hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_ready <= 1'd0;
	if (((hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_valid & (~hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_busy)) & (~hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_ready))) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_reg <= hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_payload_data;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_bitcount <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_txen & hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_busy)) begin
			hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_bitcount <= (hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_bitcount + 1'd1);
			if ((hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_busy <= 1'd0;
					hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_ready <= 1'd1;
				end else begin
					serial_tx <= hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_reg[0];
					hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_reg <= {1'd0, hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_busy) begin
		{hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_txen, hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_tx} <= (hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_tx + hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage);
	end else begin
		{hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_txen, hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_valid <= 1'd0;
	hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_r <= hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx;
	if ((~hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_busy)) begin
		if (((~hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx) & hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_r)) begin
			hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_busy <= 1'd1;
			hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_rxen) begin
			hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_bitcount <= (hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_bitcount + 1'd1);
			if ((hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_bitcount == 1'd0)) begin
				if (hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx) begin
					hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_bitcount == 4'd9)) begin
					hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_busy <= 1'd0;
					if (hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx) begin
						hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_payload_data <= hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_reg;
						hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_valid <= 1'd1;
					end
				end else begin
					hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_reg <= {hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx, hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_busy) begin
		{hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_rxen, hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_rx} <= (hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_rx + hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage);
	end else begin
		{hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_rxen, hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if (hdmi2usbsoc_hdmi2usbsoc_uart_tx_clear) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_pending <= 1'd0;
	end
	hdmi2usbsoc_hdmi2usbsoc_uart_tx_old_trigger <= hdmi2usbsoc_hdmi2usbsoc_uart_tx_trigger;
	if (((~hdmi2usbsoc_hdmi2usbsoc_uart_tx_trigger) & hdmi2usbsoc_hdmi2usbsoc_uart_tx_old_trigger)) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_pending <= 1'd1;
	end
	if (hdmi2usbsoc_hdmi2usbsoc_uart_rx_clear) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_pending <= 1'd0;
	end
	hdmi2usbsoc_hdmi2usbsoc_uart_rx_old_trigger <= hdmi2usbsoc_hdmi2usbsoc_uart_rx_trigger;
	if (((~hdmi2usbsoc_hdmi2usbsoc_uart_rx_trigger) & hdmi2usbsoc_hdmi2usbsoc_uart_rx_old_trigger)) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_pending <= 1'd1;
	end
	if (((hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_we & hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_replace))) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_produce <= (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_do_read) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_consume <= (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_we & hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_do_read)) begin
			hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level <= (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_do_read) begin
			hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level <= (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level - 1'd1);
		end
	end
	if (((hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_we & hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_replace))) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_produce <= (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_do_read) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_consume <= (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_we & hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_do_read)) begin
			hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level <= (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_do_read) begin
			hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level <= (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage) begin
		if ((hdmi2usbsoc_hdmi2usbsoc_timer0_value == 1'd0)) begin
			hdmi2usbsoc_hdmi2usbsoc_timer0_value <= hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage;
		end else begin
			hdmi2usbsoc_hdmi2usbsoc_timer0_value <= (hdmi2usbsoc_hdmi2usbsoc_timer0_value - 1'd1);
		end
	end else begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_value <= hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage;
	end
	if (hdmi2usbsoc_hdmi2usbsoc_timer0_update_value_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_value_status <= hdmi2usbsoc_hdmi2usbsoc_timer0_value;
	end
	if (hdmi2usbsoc_hdmi2usbsoc_timer0_zero_clear) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_zero_pending <= 1'd0;
	end
	hdmi2usbsoc_hdmi2usbsoc_timer0_zero_old_trigger <= hdmi2usbsoc_hdmi2usbsoc_timer0_zero_trigger;
	if (((~hdmi2usbsoc_hdmi2usbsoc_timer0_zero_trigger) & hdmi2usbsoc_hdmi2usbsoc_timer0_zero_old_trigger)) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_zero_pending <= 1'd1;
	end
	if ((hdmi2usbsoc_dna_cnt < 7'd114)) begin
		hdmi2usbsoc_dna_cnt <= (hdmi2usbsoc_dna_cnt + 1'd1);
		if (hdmi2usbsoc_dna_cnt[0]) begin
			hdmi2usbsoc_dna_status <= {hdmi2usbsoc_dna_status, hdmi2usbsoc_dna_do};
		end
	end
	if ((hdmi2usbsoc_i1 == 1'd1)) begin
		hdmi2usbsoc_clk <= 1'd1;
		hdmi2usbsoc_dqi <= hdmi2usbsoc_i0;
	end
	if ((hdmi2usbsoc_i1 == 2'd3)) begin
		hdmi2usbsoc_i1 <= 1'd0;
		hdmi2usbsoc_clk <= 1'd0;
		hdmi2usbsoc_sr <= {hdmi2usbsoc_sr[27:0], hdmi2usbsoc_dqi};
	end else begin
		hdmi2usbsoc_i1 <= (hdmi2usbsoc_i1 + 1'd1);
	end
	if ((((hdmi2usbsoc_bus_cyc & hdmi2usbsoc_bus_stb) & (hdmi2usbsoc_i1 == 2'd3)) & (hdmi2usbsoc_counter == 1'd0))) begin
		hdmi2usbsoc_dq_oe <= 1'd1;
		hdmi2usbsoc_cs_n <= 1'd0;
		hdmi2usbsoc_sr[31:0] <= 32'd4294901503;
	end
	if ((hdmi2usbsoc_counter == 6'd32)) begin
		hdmi2usbsoc_sr[31:8] <= {hdmi2usbsoc_bus_adr, {2{1'd0}}};
	end
	if ((hdmi2usbsoc_counter == 6'd56)) begin
		hdmi2usbsoc_dq_oe <= 1'd0;
	end
	if ((hdmi2usbsoc_counter == 8'd128)) begin
		hdmi2usbsoc_bus_ack <= 1'd1;
		hdmi2usbsoc_cs_n <= 1'd1;
	end
	if ((hdmi2usbsoc_counter == 8'd129)) begin
		hdmi2usbsoc_bus_ack <= 1'd0;
	end
	if ((hdmi2usbsoc_counter == 8'd133)) begin
	end
	if ((hdmi2usbsoc_counter == 8'd133)) begin
		hdmi2usbsoc_counter <= 1'd0;
	end else begin
		if ((hdmi2usbsoc_counter != 1'd0)) begin
			hdmi2usbsoc_counter <= (hdmi2usbsoc_counter + 1'd1);
		end else begin
			if (((hdmi2usbsoc_bus_cyc & hdmi2usbsoc_bus_stb) & (hdmi2usbsoc_i1 == 2'd3))) begin
				hdmi2usbsoc_counter <= 1'd1;
			end
		end
	end
	hdmi2usbsoc_ddrphy_phase_sys <= hdmi2usbsoc_ddrphy_phase_half;
	if ((hdmi2usbsoc_ddrphy_bitslip_cnt == 1'd0)) begin
		hdmi2usbsoc_ddrphy_bitslip_inc <= 1'd0;
	end else begin
		hdmi2usbsoc_ddrphy_bitslip_cnt <= (hdmi2usbsoc_ddrphy_bitslip_cnt + 1'd1);
		hdmi2usbsoc_ddrphy_bitslip_inc <= 1'd1;
	end
	hdmi2usbsoc_ddrphy_record2_wrdata <= hdmi2usbsoc_ddrphy_dfi_p0_wrdata;
	hdmi2usbsoc_ddrphy_record2_wrdata_mask <= hdmi2usbsoc_ddrphy_dfi_p0_wrdata_mask;
	hdmi2usbsoc_ddrphy_record3_wrdata <= hdmi2usbsoc_ddrphy_dfi_p1_wrdata;
	hdmi2usbsoc_ddrphy_record3_wrdata_mask <= hdmi2usbsoc_ddrphy_dfi_p1_wrdata_mask;
	hdmi2usbsoc_ddrphy_drive_dq_n1 <= hdmi2usbsoc_ddrphy_drive_dq_n0;
	hdmi2usbsoc_ddrphy_wrdata_en_d <= hdmi2usbsoc_ddrphy_wrdata_en;
	hdmi2usbsoc_ddrphy_rddata_sr <= {hdmi2usbsoc_ddrphy_rddata_en, hdmi2usbsoc_ddrphy_rddata_sr[4:1]};
	if (hdmi2usbsoc_sdram_inti_p0_rddata_valid) begin
		hdmi2usbsoc_sdram_phaseinjector0_status <= hdmi2usbsoc_sdram_inti_p0_rddata;
	end
	if (hdmi2usbsoc_sdram_inti_p1_rddata_valid) begin
		hdmi2usbsoc_sdram_phaseinjector1_status <= hdmi2usbsoc_sdram_inti_p1_rddata;
	end
	hdmi2usbsoc_sdram_cmd_payload_a <= 11'd1024;
	hdmi2usbsoc_sdram_cmd_payload_ba <= 1'd0;
	hdmi2usbsoc_sdram_cmd_payload_cas <= 1'd0;
	hdmi2usbsoc_sdram_cmd_payload_ras <= 1'd0;
	hdmi2usbsoc_sdram_cmd_payload_we <= 1'd0;
	hdmi2usbsoc_sdram_seq_done <= 1'd0;
	if ((hdmi2usbsoc_sdram_counter == 1'd1)) begin
		hdmi2usbsoc_sdram_cmd_payload_ras <= 1'd1;
		hdmi2usbsoc_sdram_cmd_payload_we <= 1'd1;
	end
	if ((hdmi2usbsoc_sdram_counter == 2'd3)) begin
		hdmi2usbsoc_sdram_cmd_payload_cas <= 1'd1;
		hdmi2usbsoc_sdram_cmd_payload_ras <= 1'd1;
	end
	if ((hdmi2usbsoc_sdram_counter == 4'd14)) begin
		hdmi2usbsoc_sdram_seq_done <= 1'd1;
	end
	if ((hdmi2usbsoc_sdram_counter == 4'd14)) begin
		hdmi2usbsoc_sdram_counter <= 1'd0;
	end else begin
		if ((hdmi2usbsoc_sdram_counter != 1'd0)) begin
			hdmi2usbsoc_sdram_counter <= (hdmi2usbsoc_sdram_counter + 1'd1);
		end else begin
			if (hdmi2usbsoc_sdram_seq_start) begin
				hdmi2usbsoc_sdram_counter <= 1'd1;
			end
		end
	end
	if (hdmi2usbsoc_sdram_wait) begin
		if ((~hdmi2usbsoc_sdram_done)) begin
			hdmi2usbsoc_sdram_count <= (hdmi2usbsoc_sdram_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_count <= 10'd585;
	end
	controllerinjector_refresher_state <= controllerinjector_refresher_next_state;
	if (hdmi2usbsoc_sdram_bankmachine0_track_close) begin
		hdmi2usbsoc_sdram_bankmachine0_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine0_track_open) begin
			hdmi2usbsoc_sdram_bankmachine0_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine0_openrow <= hdmi2usbsoc_sdram_bankmachine0_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine0_syncfifo0_we & hdmi2usbsoc_sdram_bankmachine0_syncfifo0_writable) & (~hdmi2usbsoc_sdram_bankmachine0_replace))) begin
		hdmi2usbsoc_sdram_bankmachine0_produce <= (hdmi2usbsoc_sdram_bankmachine0_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine0_do_read) begin
		hdmi2usbsoc_sdram_bankmachine0_consume <= (hdmi2usbsoc_sdram_bankmachine0_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine0_syncfifo0_we & hdmi2usbsoc_sdram_bankmachine0_syncfifo0_writable) & (~hdmi2usbsoc_sdram_bankmachine0_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine0_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine0_level <= (hdmi2usbsoc_sdram_bankmachine0_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine0_do_read) begin
			hdmi2usbsoc_sdram_bankmachine0_level <= (hdmi2usbsoc_sdram_bankmachine0_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine0_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine0_done)) begin
			hdmi2usbsoc_sdram_bankmachine0_count <= (hdmi2usbsoc_sdram_bankmachine0_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine0_count <= 3'd4;
	end
	controllerinjector_bankmachine0_state <= controllerinjector_bankmachine0_next_state;
	if (hdmi2usbsoc_sdram_bankmachine1_track_close) begin
		hdmi2usbsoc_sdram_bankmachine1_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine1_track_open) begin
			hdmi2usbsoc_sdram_bankmachine1_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine1_openrow <= hdmi2usbsoc_sdram_bankmachine1_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine1_syncfifo1_we & hdmi2usbsoc_sdram_bankmachine1_syncfifo1_writable) & (~hdmi2usbsoc_sdram_bankmachine1_replace))) begin
		hdmi2usbsoc_sdram_bankmachine1_produce <= (hdmi2usbsoc_sdram_bankmachine1_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine1_do_read) begin
		hdmi2usbsoc_sdram_bankmachine1_consume <= (hdmi2usbsoc_sdram_bankmachine1_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine1_syncfifo1_we & hdmi2usbsoc_sdram_bankmachine1_syncfifo1_writable) & (~hdmi2usbsoc_sdram_bankmachine1_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine1_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine1_level <= (hdmi2usbsoc_sdram_bankmachine1_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine1_do_read) begin
			hdmi2usbsoc_sdram_bankmachine1_level <= (hdmi2usbsoc_sdram_bankmachine1_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine1_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine1_done)) begin
			hdmi2usbsoc_sdram_bankmachine1_count <= (hdmi2usbsoc_sdram_bankmachine1_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine1_count <= 3'd4;
	end
	controllerinjector_bankmachine1_state <= controllerinjector_bankmachine1_next_state;
	if (hdmi2usbsoc_sdram_bankmachine2_track_close) begin
		hdmi2usbsoc_sdram_bankmachine2_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine2_track_open) begin
			hdmi2usbsoc_sdram_bankmachine2_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine2_openrow <= hdmi2usbsoc_sdram_bankmachine2_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine2_syncfifo2_we & hdmi2usbsoc_sdram_bankmachine2_syncfifo2_writable) & (~hdmi2usbsoc_sdram_bankmachine2_replace))) begin
		hdmi2usbsoc_sdram_bankmachine2_produce <= (hdmi2usbsoc_sdram_bankmachine2_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine2_do_read) begin
		hdmi2usbsoc_sdram_bankmachine2_consume <= (hdmi2usbsoc_sdram_bankmachine2_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine2_syncfifo2_we & hdmi2usbsoc_sdram_bankmachine2_syncfifo2_writable) & (~hdmi2usbsoc_sdram_bankmachine2_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine2_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine2_level <= (hdmi2usbsoc_sdram_bankmachine2_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine2_do_read) begin
			hdmi2usbsoc_sdram_bankmachine2_level <= (hdmi2usbsoc_sdram_bankmachine2_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine2_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine2_done)) begin
			hdmi2usbsoc_sdram_bankmachine2_count <= (hdmi2usbsoc_sdram_bankmachine2_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine2_count <= 3'd4;
	end
	controllerinjector_bankmachine2_state <= controllerinjector_bankmachine2_next_state;
	if (hdmi2usbsoc_sdram_bankmachine3_track_close) begin
		hdmi2usbsoc_sdram_bankmachine3_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine3_track_open) begin
			hdmi2usbsoc_sdram_bankmachine3_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine3_openrow <= hdmi2usbsoc_sdram_bankmachine3_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine3_syncfifo3_we & hdmi2usbsoc_sdram_bankmachine3_syncfifo3_writable) & (~hdmi2usbsoc_sdram_bankmachine3_replace))) begin
		hdmi2usbsoc_sdram_bankmachine3_produce <= (hdmi2usbsoc_sdram_bankmachine3_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine3_do_read) begin
		hdmi2usbsoc_sdram_bankmachine3_consume <= (hdmi2usbsoc_sdram_bankmachine3_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine3_syncfifo3_we & hdmi2usbsoc_sdram_bankmachine3_syncfifo3_writable) & (~hdmi2usbsoc_sdram_bankmachine3_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine3_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine3_level <= (hdmi2usbsoc_sdram_bankmachine3_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine3_do_read) begin
			hdmi2usbsoc_sdram_bankmachine3_level <= (hdmi2usbsoc_sdram_bankmachine3_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine3_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine3_done)) begin
			hdmi2usbsoc_sdram_bankmachine3_count <= (hdmi2usbsoc_sdram_bankmachine3_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine3_count <= 3'd4;
	end
	controllerinjector_bankmachine3_state <= controllerinjector_bankmachine3_next_state;
	if (hdmi2usbsoc_sdram_bankmachine4_track_close) begin
		hdmi2usbsoc_sdram_bankmachine4_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine4_track_open) begin
			hdmi2usbsoc_sdram_bankmachine4_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine4_openrow <= hdmi2usbsoc_sdram_bankmachine4_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine4_syncfifo4_we & hdmi2usbsoc_sdram_bankmachine4_syncfifo4_writable) & (~hdmi2usbsoc_sdram_bankmachine4_replace))) begin
		hdmi2usbsoc_sdram_bankmachine4_produce <= (hdmi2usbsoc_sdram_bankmachine4_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine4_do_read) begin
		hdmi2usbsoc_sdram_bankmachine4_consume <= (hdmi2usbsoc_sdram_bankmachine4_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine4_syncfifo4_we & hdmi2usbsoc_sdram_bankmachine4_syncfifo4_writable) & (~hdmi2usbsoc_sdram_bankmachine4_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine4_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine4_level <= (hdmi2usbsoc_sdram_bankmachine4_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine4_do_read) begin
			hdmi2usbsoc_sdram_bankmachine4_level <= (hdmi2usbsoc_sdram_bankmachine4_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine4_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine4_done)) begin
			hdmi2usbsoc_sdram_bankmachine4_count <= (hdmi2usbsoc_sdram_bankmachine4_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine4_count <= 3'd4;
	end
	controllerinjector_bankmachine4_state <= controllerinjector_bankmachine4_next_state;
	if (hdmi2usbsoc_sdram_bankmachine5_track_close) begin
		hdmi2usbsoc_sdram_bankmachine5_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine5_track_open) begin
			hdmi2usbsoc_sdram_bankmachine5_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine5_openrow <= hdmi2usbsoc_sdram_bankmachine5_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine5_syncfifo5_we & hdmi2usbsoc_sdram_bankmachine5_syncfifo5_writable) & (~hdmi2usbsoc_sdram_bankmachine5_replace))) begin
		hdmi2usbsoc_sdram_bankmachine5_produce <= (hdmi2usbsoc_sdram_bankmachine5_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine5_do_read) begin
		hdmi2usbsoc_sdram_bankmachine5_consume <= (hdmi2usbsoc_sdram_bankmachine5_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine5_syncfifo5_we & hdmi2usbsoc_sdram_bankmachine5_syncfifo5_writable) & (~hdmi2usbsoc_sdram_bankmachine5_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine5_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine5_level <= (hdmi2usbsoc_sdram_bankmachine5_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine5_do_read) begin
			hdmi2usbsoc_sdram_bankmachine5_level <= (hdmi2usbsoc_sdram_bankmachine5_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine5_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine5_done)) begin
			hdmi2usbsoc_sdram_bankmachine5_count <= (hdmi2usbsoc_sdram_bankmachine5_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine5_count <= 3'd4;
	end
	controllerinjector_bankmachine5_state <= controllerinjector_bankmachine5_next_state;
	if (hdmi2usbsoc_sdram_bankmachine6_track_close) begin
		hdmi2usbsoc_sdram_bankmachine6_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine6_track_open) begin
			hdmi2usbsoc_sdram_bankmachine6_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine6_openrow <= hdmi2usbsoc_sdram_bankmachine6_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine6_syncfifo6_we & hdmi2usbsoc_sdram_bankmachine6_syncfifo6_writable) & (~hdmi2usbsoc_sdram_bankmachine6_replace))) begin
		hdmi2usbsoc_sdram_bankmachine6_produce <= (hdmi2usbsoc_sdram_bankmachine6_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine6_do_read) begin
		hdmi2usbsoc_sdram_bankmachine6_consume <= (hdmi2usbsoc_sdram_bankmachine6_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine6_syncfifo6_we & hdmi2usbsoc_sdram_bankmachine6_syncfifo6_writable) & (~hdmi2usbsoc_sdram_bankmachine6_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine6_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine6_level <= (hdmi2usbsoc_sdram_bankmachine6_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine6_do_read) begin
			hdmi2usbsoc_sdram_bankmachine6_level <= (hdmi2usbsoc_sdram_bankmachine6_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine6_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine6_done)) begin
			hdmi2usbsoc_sdram_bankmachine6_count <= (hdmi2usbsoc_sdram_bankmachine6_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine6_count <= 3'd4;
	end
	controllerinjector_bankmachine6_state <= controllerinjector_bankmachine6_next_state;
	if (hdmi2usbsoc_sdram_bankmachine7_track_close) begin
		hdmi2usbsoc_sdram_bankmachine7_has_openrow <= 1'd0;
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine7_track_open) begin
			hdmi2usbsoc_sdram_bankmachine7_has_openrow <= 1'd1;
			hdmi2usbsoc_sdram_bankmachine7_openrow <= hdmi2usbsoc_sdram_bankmachine7_source_payload_adr[20:8];
		end
	end
	if (((hdmi2usbsoc_sdram_bankmachine7_syncfifo7_we & hdmi2usbsoc_sdram_bankmachine7_syncfifo7_writable) & (~hdmi2usbsoc_sdram_bankmachine7_replace))) begin
		hdmi2usbsoc_sdram_bankmachine7_produce <= (hdmi2usbsoc_sdram_bankmachine7_produce + 1'd1);
	end
	if (hdmi2usbsoc_sdram_bankmachine7_do_read) begin
		hdmi2usbsoc_sdram_bankmachine7_consume <= (hdmi2usbsoc_sdram_bankmachine7_consume + 1'd1);
	end
	if (((hdmi2usbsoc_sdram_bankmachine7_syncfifo7_we & hdmi2usbsoc_sdram_bankmachine7_syncfifo7_writable) & (~hdmi2usbsoc_sdram_bankmachine7_replace))) begin
		if ((~hdmi2usbsoc_sdram_bankmachine7_do_read)) begin
			hdmi2usbsoc_sdram_bankmachine7_level <= (hdmi2usbsoc_sdram_bankmachine7_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_sdram_bankmachine7_do_read) begin
			hdmi2usbsoc_sdram_bankmachine7_level <= (hdmi2usbsoc_sdram_bankmachine7_level - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_bankmachine7_wait) begin
		if ((~hdmi2usbsoc_sdram_bankmachine7_done)) begin
			hdmi2usbsoc_sdram_bankmachine7_count <= (hdmi2usbsoc_sdram_bankmachine7_count - 1'd1);
		end
	end else begin
		hdmi2usbsoc_sdram_bankmachine7_count <= 3'd4;
	end
	controllerinjector_bankmachine7_state <= controllerinjector_bankmachine7_next_state;
	if ((~hdmi2usbsoc_sdram_en0)) begin
		hdmi2usbsoc_sdram_time0 <= 5'd31;
	end else begin
		if ((~hdmi2usbsoc_sdram_max_time0)) begin
			hdmi2usbsoc_sdram_time0 <= (hdmi2usbsoc_sdram_time0 - 1'd1);
		end
	end
	if ((~hdmi2usbsoc_sdram_en1)) begin
		hdmi2usbsoc_sdram_time1 <= 4'd15;
	end else begin
		if ((~hdmi2usbsoc_sdram_max_time1)) begin
			hdmi2usbsoc_sdram_time1 <= (hdmi2usbsoc_sdram_time1 - 1'd1);
		end
	end
	if (hdmi2usbsoc_sdram_choose_cmd_ce) begin
		case (hdmi2usbsoc_sdram_choose_cmd_grant)
			1'd0: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[1]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd1;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[2]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd2;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[3]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd3;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[4]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd4;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[5]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd5;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[6]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd6;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[7]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[2]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd2;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[3]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd3;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[4]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd4;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[5]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd5;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[6]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd6;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[7]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd7;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[0]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[3]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd3;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[4]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd4;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[5]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd5;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[6]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd6;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[7]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd7;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[0]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd0;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[1]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[4]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd4;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[5]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd5;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[6]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd6;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[7]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd7;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[0]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd0;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[1]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd1;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[2]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[5]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd5;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[6]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd6;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[7]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd7;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[0]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd0;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[1]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd1;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[2]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd2;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[3]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[6]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd6;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[7]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd7;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[0]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd0;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[1]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd1;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[2]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd2;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[3]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd3;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[4]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[7]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd7;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[0]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd0;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[1]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd1;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[2]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd2;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[3]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd3;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[4]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd4;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[5]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (hdmi2usbsoc_sdram_choose_cmd_request[0]) begin
					hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd0;
				end else begin
					if (hdmi2usbsoc_sdram_choose_cmd_request[1]) begin
						hdmi2usbsoc_sdram_choose_cmd_grant <= 1'd1;
					end else begin
						if (hdmi2usbsoc_sdram_choose_cmd_request[2]) begin
							hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd2;
						end else begin
							if (hdmi2usbsoc_sdram_choose_cmd_request[3]) begin
								hdmi2usbsoc_sdram_choose_cmd_grant <= 2'd3;
							end else begin
								if (hdmi2usbsoc_sdram_choose_cmd_request[4]) begin
									hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd4;
								end else begin
									if (hdmi2usbsoc_sdram_choose_cmd_request[5]) begin
										hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd5;
									end else begin
										if (hdmi2usbsoc_sdram_choose_cmd_request[6]) begin
											hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (hdmi2usbsoc_sdram_choose_req_ce) begin
		case (hdmi2usbsoc_sdram_choose_req_grant)
			1'd0: begin
				if (hdmi2usbsoc_sdram_choose_req_request[1]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 1'd1;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[2]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 2'd2;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[3]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 2'd3;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[4]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 3'd4;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[5]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 3'd5;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[6]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 3'd6;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[7]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (hdmi2usbsoc_sdram_choose_req_request[2]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 2'd2;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[3]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 2'd3;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[4]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 3'd4;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[5]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 3'd5;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[6]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 3'd6;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[7]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 3'd7;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[0]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (hdmi2usbsoc_sdram_choose_req_request[3]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 2'd3;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[4]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 3'd4;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[5]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 3'd5;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[6]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 3'd6;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[7]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 3'd7;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[0]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 1'd0;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[1]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (hdmi2usbsoc_sdram_choose_req_request[4]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 3'd4;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[5]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 3'd5;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[6]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 3'd6;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[7]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 3'd7;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[0]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 1'd0;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[1]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 1'd1;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[2]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (hdmi2usbsoc_sdram_choose_req_request[5]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 3'd5;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[6]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 3'd6;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[7]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 3'd7;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[0]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 1'd0;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[1]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 1'd1;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[2]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 2'd2;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[3]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (hdmi2usbsoc_sdram_choose_req_request[6]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 3'd6;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[7]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 3'd7;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[0]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 1'd0;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[1]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 1'd1;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[2]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 2'd2;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[3]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 2'd3;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[4]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (hdmi2usbsoc_sdram_choose_req_request[7]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 3'd7;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[0]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 1'd0;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[1]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 1'd1;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[2]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 2'd2;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[3]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 2'd3;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[4]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 3'd4;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[5]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (hdmi2usbsoc_sdram_choose_req_request[0]) begin
					hdmi2usbsoc_sdram_choose_req_grant <= 1'd0;
				end else begin
					if (hdmi2usbsoc_sdram_choose_req_request[1]) begin
						hdmi2usbsoc_sdram_choose_req_grant <= 1'd1;
					end else begin
						if (hdmi2usbsoc_sdram_choose_req_request[2]) begin
							hdmi2usbsoc_sdram_choose_req_grant <= 2'd2;
						end else begin
							if (hdmi2usbsoc_sdram_choose_req_request[3]) begin
								hdmi2usbsoc_sdram_choose_req_grant <= 2'd3;
							end else begin
								if (hdmi2usbsoc_sdram_choose_req_request[4]) begin
									hdmi2usbsoc_sdram_choose_req_grant <= 3'd4;
								end else begin
									if (hdmi2usbsoc_sdram_choose_req_request[5]) begin
										hdmi2usbsoc_sdram_choose_req_grant <= 3'd5;
									end else begin
										if (hdmi2usbsoc_sdram_choose_req_request[6]) begin
											hdmi2usbsoc_sdram_choose_req_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	hdmi2usbsoc_sdram_dfi_p0_address <= sync_rhs_array_muxed7;
	hdmi2usbsoc_sdram_dfi_p0_bank <= sync_rhs_array_muxed8;
	hdmi2usbsoc_sdram_dfi_p0_cas_n <= (~sync_rhs_array_muxed9);
	hdmi2usbsoc_sdram_dfi_p0_ras_n <= (~sync_rhs_array_muxed10);
	hdmi2usbsoc_sdram_dfi_p0_we_n <= (~sync_rhs_array_muxed11);
	hdmi2usbsoc_sdram_dfi_p0_rddata_en <= sync_rhs_array_muxed12;
	hdmi2usbsoc_sdram_dfi_p0_wrdata_en <= sync_rhs_array_muxed13;
	hdmi2usbsoc_sdram_dfi_p1_address <= sync_rhs_array_muxed14;
	hdmi2usbsoc_sdram_dfi_p1_bank <= sync_rhs_array_muxed15;
	hdmi2usbsoc_sdram_dfi_p1_cas_n <= (~sync_rhs_array_muxed16);
	hdmi2usbsoc_sdram_dfi_p1_ras_n <= (~sync_rhs_array_muxed17);
	hdmi2usbsoc_sdram_dfi_p1_we_n <= (~sync_rhs_array_muxed18);
	hdmi2usbsoc_sdram_dfi_p1_rddata_en <= sync_rhs_array_muxed19;
	hdmi2usbsoc_sdram_dfi_p1_wrdata_en <= sync_rhs_array_muxed20;
	controllerinjector_multiplexer_state <= controllerinjector_multiplexer_next_state;
	hdmi2usbsoc_sdram_bandwidth_cmd_valid <= hdmi2usbsoc_sdram_choose_req_cmd_valid;
	hdmi2usbsoc_sdram_bandwidth_cmd_ready <= hdmi2usbsoc_sdram_choose_req_cmd_ready;
	hdmi2usbsoc_sdram_bandwidth_cmd_is_read <= hdmi2usbsoc_sdram_choose_req_cmd_payload_is_read;
	hdmi2usbsoc_sdram_bandwidth_cmd_is_write <= hdmi2usbsoc_sdram_choose_req_cmd_payload_is_write;
	{hdmi2usbsoc_sdram_bandwidth_period, hdmi2usbsoc_sdram_bandwidth_counter} <= (hdmi2usbsoc_sdram_bandwidth_counter + 1'd1);
	if (hdmi2usbsoc_sdram_bandwidth_period) begin
		hdmi2usbsoc_sdram_bandwidth_nreads_r <= hdmi2usbsoc_sdram_bandwidth_nreads;
		hdmi2usbsoc_sdram_bandwidth_nwrites_r <= hdmi2usbsoc_sdram_bandwidth_nwrites;
		hdmi2usbsoc_sdram_bandwidth_nreads <= 1'd0;
		hdmi2usbsoc_sdram_bandwidth_nwrites <= 1'd0;
	end else begin
		if ((hdmi2usbsoc_sdram_bandwidth_cmd_valid & hdmi2usbsoc_sdram_bandwidth_cmd_ready)) begin
			if (hdmi2usbsoc_sdram_bandwidth_cmd_is_read) begin
				hdmi2usbsoc_sdram_bandwidth_nreads <= (hdmi2usbsoc_sdram_bandwidth_nreads + 1'd1);
			end
			if (hdmi2usbsoc_sdram_bandwidth_cmd_is_write) begin
				hdmi2usbsoc_sdram_bandwidth_nwrites <= (hdmi2usbsoc_sdram_bandwidth_nwrites + 1'd1);
			end
		end
	end
	if (hdmi2usbsoc_sdram_bandwidth_update_re) begin
		hdmi2usbsoc_sdram_bandwidth_nreads_status <= hdmi2usbsoc_sdram_bandwidth_nreads_r;
		hdmi2usbsoc_sdram_bandwidth_nwrites_status <= hdmi2usbsoc_sdram_bandwidth_nwrites_r;
	end
	controllerinjector_new_master_wdata_ready0 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank0_wdata_ready)) | ((controllerinjector_roundrobin1_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank1_wdata_ready)) | ((controllerinjector_roundrobin2_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank2_wdata_ready)) | ((controllerinjector_roundrobin3_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank3_wdata_ready)) | ((controllerinjector_roundrobin4_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank4_wdata_ready)) | ((controllerinjector_roundrobin5_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank5_wdata_ready)) | ((controllerinjector_roundrobin6_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank6_wdata_ready)) | ((controllerinjector_roundrobin7_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank7_wdata_ready));
	controllerinjector_new_master_wdata_ready1 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank0_wdata_ready)) | ((controllerinjector_roundrobin1_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank1_wdata_ready)) | ((controllerinjector_roundrobin2_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank2_wdata_ready)) | ((controllerinjector_roundrobin3_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank3_wdata_ready)) | ((controllerinjector_roundrobin4_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank4_wdata_ready)) | ((controllerinjector_roundrobin5_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank5_wdata_ready)) | ((controllerinjector_roundrobin6_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank6_wdata_ready)) | ((controllerinjector_roundrobin7_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank7_wdata_ready));
	controllerinjector_new_master_wdata_ready2 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank0_wdata_ready)) | ((controllerinjector_roundrobin1_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank1_wdata_ready)) | ((controllerinjector_roundrobin2_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank2_wdata_ready)) | ((controllerinjector_roundrobin3_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank3_wdata_ready)) | ((controllerinjector_roundrobin4_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank4_wdata_ready)) | ((controllerinjector_roundrobin5_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank5_wdata_ready)) | ((controllerinjector_roundrobin6_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank6_wdata_ready)) | ((controllerinjector_roundrobin7_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank7_wdata_ready));
	controllerinjector_new_master_wdata_ready3 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank0_wdata_ready)) | ((controllerinjector_roundrobin1_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank1_wdata_ready)) | ((controllerinjector_roundrobin2_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank2_wdata_ready)) | ((controllerinjector_roundrobin3_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank3_wdata_ready)) | ((controllerinjector_roundrobin4_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank4_wdata_ready)) | ((controllerinjector_roundrobin5_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank5_wdata_ready)) | ((controllerinjector_roundrobin6_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank6_wdata_ready)) | ((controllerinjector_roundrobin7_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank7_wdata_ready));
	controllerinjector_new_master_wdata_ready4 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank0_wdata_ready)) | ((controllerinjector_roundrobin1_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank1_wdata_ready)) | ((controllerinjector_roundrobin2_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank2_wdata_ready)) | ((controllerinjector_roundrobin3_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank3_wdata_ready)) | ((controllerinjector_roundrobin4_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank4_wdata_ready)) | ((controllerinjector_roundrobin5_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank5_wdata_ready)) | ((controllerinjector_roundrobin6_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank6_wdata_ready)) | ((controllerinjector_roundrobin7_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank7_wdata_ready));
	controllerinjector_new_master_wdata_ready5 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank0_wdata_ready)) | ((controllerinjector_roundrobin1_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank1_wdata_ready)) | ((controllerinjector_roundrobin2_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank2_wdata_ready)) | ((controllerinjector_roundrobin3_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank3_wdata_ready)) | ((controllerinjector_roundrobin4_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank4_wdata_ready)) | ((controllerinjector_roundrobin5_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank5_wdata_ready)) | ((controllerinjector_roundrobin6_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank6_wdata_ready)) | ((controllerinjector_roundrobin7_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank7_wdata_ready));
	controllerinjector_new_master_rdata_valid0 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank0_rdata_valid)) | ((controllerinjector_roundrobin1_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank1_rdata_valid)) | ((controllerinjector_roundrobin2_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank2_rdata_valid)) | ((controllerinjector_roundrobin3_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank3_rdata_valid)) | ((controllerinjector_roundrobin4_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank4_rdata_valid)) | ((controllerinjector_roundrobin5_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank5_rdata_valid)) | ((controllerinjector_roundrobin6_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank6_rdata_valid)) | ((controllerinjector_roundrobin7_grant == 1'd0) & hdmi2usbsoc_sdram_interface_bank7_rdata_valid));
	controllerinjector_new_master_rdata_valid1 <= controllerinjector_new_master_rdata_valid0;
	controllerinjector_new_master_rdata_valid2 <= controllerinjector_new_master_rdata_valid1;
	controllerinjector_new_master_rdata_valid3 <= controllerinjector_new_master_rdata_valid2;
	controllerinjector_new_master_rdata_valid4 <= controllerinjector_new_master_rdata_valid3;
	controllerinjector_new_master_rdata_valid5 <= controllerinjector_new_master_rdata_valid4;
	controllerinjector_new_master_rdata_valid6 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank0_rdata_valid)) | ((controllerinjector_roundrobin1_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank1_rdata_valid)) | ((controllerinjector_roundrobin2_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank2_rdata_valid)) | ((controllerinjector_roundrobin3_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank3_rdata_valid)) | ((controllerinjector_roundrobin4_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank4_rdata_valid)) | ((controllerinjector_roundrobin5_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank5_rdata_valid)) | ((controllerinjector_roundrobin6_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank6_rdata_valid)) | ((controllerinjector_roundrobin7_grant == 1'd1) & hdmi2usbsoc_sdram_interface_bank7_rdata_valid));
	controllerinjector_new_master_rdata_valid7 <= controllerinjector_new_master_rdata_valid6;
	controllerinjector_new_master_rdata_valid8 <= controllerinjector_new_master_rdata_valid7;
	controllerinjector_new_master_rdata_valid9 <= controllerinjector_new_master_rdata_valid8;
	controllerinjector_new_master_rdata_valid10 <= controllerinjector_new_master_rdata_valid9;
	controllerinjector_new_master_rdata_valid11 <= controllerinjector_new_master_rdata_valid10;
	controllerinjector_new_master_rdata_valid12 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank0_rdata_valid)) | ((controllerinjector_roundrobin1_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank1_rdata_valid)) | ((controllerinjector_roundrobin2_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank2_rdata_valid)) | ((controllerinjector_roundrobin3_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank3_rdata_valid)) | ((controllerinjector_roundrobin4_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank4_rdata_valid)) | ((controllerinjector_roundrobin5_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank5_rdata_valid)) | ((controllerinjector_roundrobin6_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank6_rdata_valid)) | ((controllerinjector_roundrobin7_grant == 2'd2) & hdmi2usbsoc_sdram_interface_bank7_rdata_valid));
	controllerinjector_new_master_rdata_valid13 <= controllerinjector_new_master_rdata_valid12;
	controllerinjector_new_master_rdata_valid14 <= controllerinjector_new_master_rdata_valid13;
	controllerinjector_new_master_rdata_valid15 <= controllerinjector_new_master_rdata_valid14;
	controllerinjector_new_master_rdata_valid16 <= controllerinjector_new_master_rdata_valid15;
	controllerinjector_new_master_rdata_valid17 <= controllerinjector_new_master_rdata_valid16;
	controllerinjector_new_master_rdata_valid18 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank0_rdata_valid)) | ((controllerinjector_roundrobin1_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank1_rdata_valid)) | ((controllerinjector_roundrobin2_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank2_rdata_valid)) | ((controllerinjector_roundrobin3_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank3_rdata_valid)) | ((controllerinjector_roundrobin4_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank4_rdata_valid)) | ((controllerinjector_roundrobin5_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank5_rdata_valid)) | ((controllerinjector_roundrobin6_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank6_rdata_valid)) | ((controllerinjector_roundrobin7_grant == 2'd3) & hdmi2usbsoc_sdram_interface_bank7_rdata_valid));
	controllerinjector_new_master_rdata_valid19 <= controllerinjector_new_master_rdata_valid18;
	controllerinjector_new_master_rdata_valid20 <= controllerinjector_new_master_rdata_valid19;
	controllerinjector_new_master_rdata_valid21 <= controllerinjector_new_master_rdata_valid20;
	controllerinjector_new_master_rdata_valid22 <= controllerinjector_new_master_rdata_valid21;
	controllerinjector_new_master_rdata_valid23 <= controllerinjector_new_master_rdata_valid22;
	controllerinjector_new_master_rdata_valid24 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank0_rdata_valid)) | ((controllerinjector_roundrobin1_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank1_rdata_valid)) | ((controllerinjector_roundrobin2_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank2_rdata_valid)) | ((controllerinjector_roundrobin3_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank3_rdata_valid)) | ((controllerinjector_roundrobin4_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank4_rdata_valid)) | ((controllerinjector_roundrobin5_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank5_rdata_valid)) | ((controllerinjector_roundrobin6_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank6_rdata_valid)) | ((controllerinjector_roundrobin7_grant == 3'd4) & hdmi2usbsoc_sdram_interface_bank7_rdata_valid));
	controllerinjector_new_master_rdata_valid25 <= controllerinjector_new_master_rdata_valid24;
	controllerinjector_new_master_rdata_valid26 <= controllerinjector_new_master_rdata_valid25;
	controllerinjector_new_master_rdata_valid27 <= controllerinjector_new_master_rdata_valid26;
	controllerinjector_new_master_rdata_valid28 <= controllerinjector_new_master_rdata_valid27;
	controllerinjector_new_master_rdata_valid29 <= controllerinjector_new_master_rdata_valid28;
	controllerinjector_new_master_rdata_valid30 <= ((((((((1'd0 | ((controllerinjector_roundrobin0_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank0_rdata_valid)) | ((controllerinjector_roundrobin1_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank1_rdata_valid)) | ((controllerinjector_roundrobin2_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank2_rdata_valid)) | ((controllerinjector_roundrobin3_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank3_rdata_valid)) | ((controllerinjector_roundrobin4_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank4_rdata_valid)) | ((controllerinjector_roundrobin5_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank5_rdata_valid)) | ((controllerinjector_roundrobin6_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank6_rdata_valid)) | ((controllerinjector_roundrobin7_grant == 3'd5) & hdmi2usbsoc_sdram_interface_bank7_rdata_valid));
	controllerinjector_new_master_rdata_valid31 <= controllerinjector_new_master_rdata_valid30;
	controllerinjector_new_master_rdata_valid32 <= controllerinjector_new_master_rdata_valid31;
	controllerinjector_new_master_rdata_valid33 <= controllerinjector_new_master_rdata_valid32;
	controllerinjector_new_master_rdata_valid34 <= controllerinjector_new_master_rdata_valid33;
	controllerinjector_new_master_rdata_valid35 <= controllerinjector_new_master_rdata_valid34;
	hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_binary <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next_binary;
	hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_next;
	hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_binary <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next_binary;
	hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_next;
	hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_binary <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next_binary;
	hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_next;
	hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_binary <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next_binary;
	hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_next;
	if (encoder_port_counter_reset) begin
		encoder_port_counter <= 1'd0;
	end else begin
		if (encoder_port_counter_ce) begin
			encoder_port_counter <= (encoder_port_counter + 1'd1);
		end
	end
	controllerinjector_state <= controllerinjector_next_state;
	if (encoder_port_converter_source_ready) begin
		encoder_port_converter_strobe_all <= 1'd0;
	end
	if (encoder_port_converter_load_part) begin
		if (((encoder_port_converter_demux == 1'd1) | encoder_port_converter_sink_last)) begin
			encoder_port_converter_demux <= 1'd0;
			encoder_port_converter_strobe_all <= 1'd1;
		end else begin
			encoder_port_converter_demux <= (encoder_port_converter_demux + 1'd1);
		end
	end
	if ((encoder_port_converter_source_valid & encoder_port_converter_source_ready)) begin
		if ((encoder_port_converter_sink_valid & encoder_port_converter_sink_ready)) begin
			encoder_port_converter_source_first <= encoder_port_converter_sink_first;
			encoder_port_converter_source_last <= encoder_port_converter_sink_last;
		end else begin
			encoder_port_converter_source_first <= 1'd0;
			encoder_port_converter_source_last <= 1'd0;
		end
	end else begin
		if ((encoder_port_converter_sink_valid & encoder_port_converter_sink_ready)) begin
			encoder_port_converter_source_first <= (encoder_port_converter_sink_first | encoder_port_converter_source_first);
			encoder_port_converter_source_last <= (encoder_port_converter_sink_last | encoder_port_converter_source_last);
		end
	end
	if (encoder_port_converter_load_part) begin
		case (encoder_port_converter_demux)
			1'd0: begin
				encoder_port_converter_source_payload_data[127:64] <= encoder_port_converter_sink_payload_data;
			end
			1'd1: begin
				encoder_port_converter_source_payload_data[63:0] <= encoder_port_converter_sink_payload_data;
			end
		endcase
	end
	if (encoder_port_converter_load_part) begin
		encoder_port_converter_source_payload_valid_token_count <= (encoder_port_converter_demux + 1'd1);
	end
	if (controllerinjector_roundrobin0_ce) begin
		case (controllerinjector_roundrobin0_grant)
			1'd0: begin
				if (controllerinjector_roundrobin0_request[1]) begin
					controllerinjector_roundrobin0_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin0_request[2]) begin
						controllerinjector_roundrobin0_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin0_request[3]) begin
							controllerinjector_roundrobin0_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin0_request[4]) begin
								controllerinjector_roundrobin0_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin0_request[5]) begin
									controllerinjector_roundrobin0_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin0_request[2]) begin
					controllerinjector_roundrobin0_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin0_request[3]) begin
						controllerinjector_roundrobin0_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin0_request[4]) begin
							controllerinjector_roundrobin0_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin0_request[5]) begin
								controllerinjector_roundrobin0_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin0_request[0]) begin
									controllerinjector_roundrobin0_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin0_request[3]) begin
					controllerinjector_roundrobin0_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin0_request[4]) begin
						controllerinjector_roundrobin0_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin0_request[5]) begin
							controllerinjector_roundrobin0_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin0_request[0]) begin
								controllerinjector_roundrobin0_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin0_request[1]) begin
									controllerinjector_roundrobin0_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin0_request[4]) begin
					controllerinjector_roundrobin0_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin0_request[5]) begin
						controllerinjector_roundrobin0_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin0_request[0]) begin
							controllerinjector_roundrobin0_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin0_request[1]) begin
								controllerinjector_roundrobin0_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin0_request[2]) begin
									controllerinjector_roundrobin0_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin0_request[5]) begin
					controllerinjector_roundrobin0_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin0_request[0]) begin
						controllerinjector_roundrobin0_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin0_request[1]) begin
							controllerinjector_roundrobin0_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin0_request[2]) begin
								controllerinjector_roundrobin0_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin0_request[3]) begin
									controllerinjector_roundrobin0_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin0_request[0]) begin
					controllerinjector_roundrobin0_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin0_request[1]) begin
						controllerinjector_roundrobin0_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin0_request[2]) begin
							controllerinjector_roundrobin0_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin0_request[3]) begin
								controllerinjector_roundrobin0_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin0_request[4]) begin
									controllerinjector_roundrobin0_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (controllerinjector_roundrobin1_ce) begin
		case (controllerinjector_roundrobin1_grant)
			1'd0: begin
				if (controllerinjector_roundrobin1_request[1]) begin
					controllerinjector_roundrobin1_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin1_request[2]) begin
						controllerinjector_roundrobin1_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin1_request[3]) begin
							controllerinjector_roundrobin1_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin1_request[4]) begin
								controllerinjector_roundrobin1_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin1_request[5]) begin
									controllerinjector_roundrobin1_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin1_request[2]) begin
					controllerinjector_roundrobin1_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin1_request[3]) begin
						controllerinjector_roundrobin1_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin1_request[4]) begin
							controllerinjector_roundrobin1_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin1_request[5]) begin
								controllerinjector_roundrobin1_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin1_request[0]) begin
									controllerinjector_roundrobin1_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin1_request[3]) begin
					controllerinjector_roundrobin1_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin1_request[4]) begin
						controllerinjector_roundrobin1_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin1_request[5]) begin
							controllerinjector_roundrobin1_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin1_request[0]) begin
								controllerinjector_roundrobin1_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin1_request[1]) begin
									controllerinjector_roundrobin1_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin1_request[4]) begin
					controllerinjector_roundrobin1_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin1_request[5]) begin
						controllerinjector_roundrobin1_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin1_request[0]) begin
							controllerinjector_roundrobin1_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin1_request[1]) begin
								controllerinjector_roundrobin1_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin1_request[2]) begin
									controllerinjector_roundrobin1_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin1_request[5]) begin
					controllerinjector_roundrobin1_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin1_request[0]) begin
						controllerinjector_roundrobin1_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin1_request[1]) begin
							controllerinjector_roundrobin1_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin1_request[2]) begin
								controllerinjector_roundrobin1_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin1_request[3]) begin
									controllerinjector_roundrobin1_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin1_request[0]) begin
					controllerinjector_roundrobin1_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin1_request[1]) begin
						controllerinjector_roundrobin1_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin1_request[2]) begin
							controllerinjector_roundrobin1_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin1_request[3]) begin
								controllerinjector_roundrobin1_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin1_request[4]) begin
									controllerinjector_roundrobin1_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (controllerinjector_roundrobin2_ce) begin
		case (controllerinjector_roundrobin2_grant)
			1'd0: begin
				if (controllerinjector_roundrobin2_request[1]) begin
					controllerinjector_roundrobin2_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin2_request[2]) begin
						controllerinjector_roundrobin2_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin2_request[3]) begin
							controllerinjector_roundrobin2_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin2_request[4]) begin
								controllerinjector_roundrobin2_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin2_request[5]) begin
									controllerinjector_roundrobin2_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin2_request[2]) begin
					controllerinjector_roundrobin2_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin2_request[3]) begin
						controllerinjector_roundrobin2_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin2_request[4]) begin
							controllerinjector_roundrobin2_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin2_request[5]) begin
								controllerinjector_roundrobin2_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin2_request[0]) begin
									controllerinjector_roundrobin2_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin2_request[3]) begin
					controllerinjector_roundrobin2_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin2_request[4]) begin
						controllerinjector_roundrobin2_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin2_request[5]) begin
							controllerinjector_roundrobin2_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin2_request[0]) begin
								controllerinjector_roundrobin2_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin2_request[1]) begin
									controllerinjector_roundrobin2_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin2_request[4]) begin
					controllerinjector_roundrobin2_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin2_request[5]) begin
						controllerinjector_roundrobin2_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin2_request[0]) begin
							controllerinjector_roundrobin2_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin2_request[1]) begin
								controllerinjector_roundrobin2_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin2_request[2]) begin
									controllerinjector_roundrobin2_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin2_request[5]) begin
					controllerinjector_roundrobin2_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin2_request[0]) begin
						controllerinjector_roundrobin2_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin2_request[1]) begin
							controllerinjector_roundrobin2_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin2_request[2]) begin
								controllerinjector_roundrobin2_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin2_request[3]) begin
									controllerinjector_roundrobin2_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin2_request[0]) begin
					controllerinjector_roundrobin2_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin2_request[1]) begin
						controllerinjector_roundrobin2_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin2_request[2]) begin
							controllerinjector_roundrobin2_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin2_request[3]) begin
								controllerinjector_roundrobin2_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin2_request[4]) begin
									controllerinjector_roundrobin2_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (controllerinjector_roundrobin3_ce) begin
		case (controllerinjector_roundrobin3_grant)
			1'd0: begin
				if (controllerinjector_roundrobin3_request[1]) begin
					controllerinjector_roundrobin3_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin3_request[2]) begin
						controllerinjector_roundrobin3_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin3_request[3]) begin
							controllerinjector_roundrobin3_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin3_request[4]) begin
								controllerinjector_roundrobin3_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin3_request[5]) begin
									controllerinjector_roundrobin3_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin3_request[2]) begin
					controllerinjector_roundrobin3_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin3_request[3]) begin
						controllerinjector_roundrobin3_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin3_request[4]) begin
							controllerinjector_roundrobin3_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin3_request[5]) begin
								controllerinjector_roundrobin3_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin3_request[0]) begin
									controllerinjector_roundrobin3_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin3_request[3]) begin
					controllerinjector_roundrobin3_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin3_request[4]) begin
						controllerinjector_roundrobin3_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin3_request[5]) begin
							controllerinjector_roundrobin3_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin3_request[0]) begin
								controllerinjector_roundrobin3_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin3_request[1]) begin
									controllerinjector_roundrobin3_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin3_request[4]) begin
					controllerinjector_roundrobin3_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin3_request[5]) begin
						controllerinjector_roundrobin3_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin3_request[0]) begin
							controllerinjector_roundrobin3_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin3_request[1]) begin
								controllerinjector_roundrobin3_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin3_request[2]) begin
									controllerinjector_roundrobin3_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin3_request[5]) begin
					controllerinjector_roundrobin3_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin3_request[0]) begin
						controllerinjector_roundrobin3_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin3_request[1]) begin
							controllerinjector_roundrobin3_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin3_request[2]) begin
								controllerinjector_roundrobin3_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin3_request[3]) begin
									controllerinjector_roundrobin3_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin3_request[0]) begin
					controllerinjector_roundrobin3_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin3_request[1]) begin
						controllerinjector_roundrobin3_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin3_request[2]) begin
							controllerinjector_roundrobin3_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin3_request[3]) begin
								controllerinjector_roundrobin3_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin3_request[4]) begin
									controllerinjector_roundrobin3_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (controllerinjector_roundrobin4_ce) begin
		case (controllerinjector_roundrobin4_grant)
			1'd0: begin
				if (controllerinjector_roundrobin4_request[1]) begin
					controllerinjector_roundrobin4_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin4_request[2]) begin
						controllerinjector_roundrobin4_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin4_request[3]) begin
							controllerinjector_roundrobin4_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin4_request[4]) begin
								controllerinjector_roundrobin4_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin4_request[5]) begin
									controllerinjector_roundrobin4_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin4_request[2]) begin
					controllerinjector_roundrobin4_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin4_request[3]) begin
						controllerinjector_roundrobin4_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin4_request[4]) begin
							controllerinjector_roundrobin4_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin4_request[5]) begin
								controllerinjector_roundrobin4_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin4_request[0]) begin
									controllerinjector_roundrobin4_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin4_request[3]) begin
					controllerinjector_roundrobin4_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin4_request[4]) begin
						controllerinjector_roundrobin4_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin4_request[5]) begin
							controllerinjector_roundrobin4_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin4_request[0]) begin
								controllerinjector_roundrobin4_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin4_request[1]) begin
									controllerinjector_roundrobin4_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin4_request[4]) begin
					controllerinjector_roundrobin4_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin4_request[5]) begin
						controllerinjector_roundrobin4_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin4_request[0]) begin
							controllerinjector_roundrobin4_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin4_request[1]) begin
								controllerinjector_roundrobin4_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin4_request[2]) begin
									controllerinjector_roundrobin4_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin4_request[5]) begin
					controllerinjector_roundrobin4_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin4_request[0]) begin
						controllerinjector_roundrobin4_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin4_request[1]) begin
							controllerinjector_roundrobin4_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin4_request[2]) begin
								controllerinjector_roundrobin4_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin4_request[3]) begin
									controllerinjector_roundrobin4_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin4_request[0]) begin
					controllerinjector_roundrobin4_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin4_request[1]) begin
						controllerinjector_roundrobin4_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin4_request[2]) begin
							controllerinjector_roundrobin4_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin4_request[3]) begin
								controllerinjector_roundrobin4_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin4_request[4]) begin
									controllerinjector_roundrobin4_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (controllerinjector_roundrobin5_ce) begin
		case (controllerinjector_roundrobin5_grant)
			1'd0: begin
				if (controllerinjector_roundrobin5_request[1]) begin
					controllerinjector_roundrobin5_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin5_request[2]) begin
						controllerinjector_roundrobin5_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin5_request[3]) begin
							controllerinjector_roundrobin5_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin5_request[4]) begin
								controllerinjector_roundrobin5_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin5_request[5]) begin
									controllerinjector_roundrobin5_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin5_request[2]) begin
					controllerinjector_roundrobin5_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin5_request[3]) begin
						controllerinjector_roundrobin5_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin5_request[4]) begin
							controllerinjector_roundrobin5_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin5_request[5]) begin
								controllerinjector_roundrobin5_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin5_request[0]) begin
									controllerinjector_roundrobin5_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin5_request[3]) begin
					controllerinjector_roundrobin5_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin5_request[4]) begin
						controllerinjector_roundrobin5_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin5_request[5]) begin
							controllerinjector_roundrobin5_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin5_request[0]) begin
								controllerinjector_roundrobin5_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin5_request[1]) begin
									controllerinjector_roundrobin5_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin5_request[4]) begin
					controllerinjector_roundrobin5_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin5_request[5]) begin
						controllerinjector_roundrobin5_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin5_request[0]) begin
							controllerinjector_roundrobin5_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin5_request[1]) begin
								controllerinjector_roundrobin5_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin5_request[2]) begin
									controllerinjector_roundrobin5_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin5_request[5]) begin
					controllerinjector_roundrobin5_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin5_request[0]) begin
						controllerinjector_roundrobin5_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin5_request[1]) begin
							controllerinjector_roundrobin5_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin5_request[2]) begin
								controllerinjector_roundrobin5_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin5_request[3]) begin
									controllerinjector_roundrobin5_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin5_request[0]) begin
					controllerinjector_roundrobin5_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin5_request[1]) begin
						controllerinjector_roundrobin5_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin5_request[2]) begin
							controllerinjector_roundrobin5_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin5_request[3]) begin
								controllerinjector_roundrobin5_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin5_request[4]) begin
									controllerinjector_roundrobin5_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (controllerinjector_roundrobin6_ce) begin
		case (controllerinjector_roundrobin6_grant)
			1'd0: begin
				if (controllerinjector_roundrobin6_request[1]) begin
					controllerinjector_roundrobin6_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin6_request[2]) begin
						controllerinjector_roundrobin6_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin6_request[3]) begin
							controllerinjector_roundrobin6_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin6_request[4]) begin
								controllerinjector_roundrobin6_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin6_request[5]) begin
									controllerinjector_roundrobin6_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin6_request[2]) begin
					controllerinjector_roundrobin6_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin6_request[3]) begin
						controllerinjector_roundrobin6_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin6_request[4]) begin
							controllerinjector_roundrobin6_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin6_request[5]) begin
								controllerinjector_roundrobin6_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin6_request[0]) begin
									controllerinjector_roundrobin6_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin6_request[3]) begin
					controllerinjector_roundrobin6_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin6_request[4]) begin
						controllerinjector_roundrobin6_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin6_request[5]) begin
							controllerinjector_roundrobin6_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin6_request[0]) begin
								controllerinjector_roundrobin6_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin6_request[1]) begin
									controllerinjector_roundrobin6_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin6_request[4]) begin
					controllerinjector_roundrobin6_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin6_request[5]) begin
						controllerinjector_roundrobin6_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin6_request[0]) begin
							controllerinjector_roundrobin6_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin6_request[1]) begin
								controllerinjector_roundrobin6_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin6_request[2]) begin
									controllerinjector_roundrobin6_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin6_request[5]) begin
					controllerinjector_roundrobin6_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin6_request[0]) begin
						controllerinjector_roundrobin6_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin6_request[1]) begin
							controllerinjector_roundrobin6_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin6_request[2]) begin
								controllerinjector_roundrobin6_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin6_request[3]) begin
									controllerinjector_roundrobin6_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin6_request[0]) begin
					controllerinjector_roundrobin6_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin6_request[1]) begin
						controllerinjector_roundrobin6_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin6_request[2]) begin
							controllerinjector_roundrobin6_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin6_request[3]) begin
								controllerinjector_roundrobin6_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin6_request[4]) begin
									controllerinjector_roundrobin6_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (controllerinjector_roundrobin7_ce) begin
		case (controllerinjector_roundrobin7_grant)
			1'd0: begin
				if (controllerinjector_roundrobin7_request[1]) begin
					controllerinjector_roundrobin7_grant <= 1'd1;
				end else begin
					if (controllerinjector_roundrobin7_request[2]) begin
						controllerinjector_roundrobin7_grant <= 2'd2;
					end else begin
						if (controllerinjector_roundrobin7_request[3]) begin
							controllerinjector_roundrobin7_grant <= 2'd3;
						end else begin
							if (controllerinjector_roundrobin7_request[4]) begin
								controllerinjector_roundrobin7_grant <= 3'd4;
							end else begin
								if (controllerinjector_roundrobin7_request[5]) begin
									controllerinjector_roundrobin7_grant <= 3'd5;
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (controllerinjector_roundrobin7_request[2]) begin
					controllerinjector_roundrobin7_grant <= 2'd2;
				end else begin
					if (controllerinjector_roundrobin7_request[3]) begin
						controllerinjector_roundrobin7_grant <= 2'd3;
					end else begin
						if (controllerinjector_roundrobin7_request[4]) begin
							controllerinjector_roundrobin7_grant <= 3'd4;
						end else begin
							if (controllerinjector_roundrobin7_request[5]) begin
								controllerinjector_roundrobin7_grant <= 3'd5;
							end else begin
								if (controllerinjector_roundrobin7_request[0]) begin
									controllerinjector_roundrobin7_grant <= 1'd0;
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (controllerinjector_roundrobin7_request[3]) begin
					controllerinjector_roundrobin7_grant <= 2'd3;
				end else begin
					if (controllerinjector_roundrobin7_request[4]) begin
						controllerinjector_roundrobin7_grant <= 3'd4;
					end else begin
						if (controllerinjector_roundrobin7_request[5]) begin
							controllerinjector_roundrobin7_grant <= 3'd5;
						end else begin
							if (controllerinjector_roundrobin7_request[0]) begin
								controllerinjector_roundrobin7_grant <= 1'd0;
							end else begin
								if (controllerinjector_roundrobin7_request[1]) begin
									controllerinjector_roundrobin7_grant <= 1'd1;
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (controllerinjector_roundrobin7_request[4]) begin
					controllerinjector_roundrobin7_grant <= 3'd4;
				end else begin
					if (controllerinjector_roundrobin7_request[5]) begin
						controllerinjector_roundrobin7_grant <= 3'd5;
					end else begin
						if (controllerinjector_roundrobin7_request[0]) begin
							controllerinjector_roundrobin7_grant <= 1'd0;
						end else begin
							if (controllerinjector_roundrobin7_request[1]) begin
								controllerinjector_roundrobin7_grant <= 1'd1;
							end else begin
								if (controllerinjector_roundrobin7_request[2]) begin
									controllerinjector_roundrobin7_grant <= 2'd2;
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (controllerinjector_roundrobin7_request[5]) begin
					controllerinjector_roundrobin7_grant <= 3'd5;
				end else begin
					if (controllerinjector_roundrobin7_request[0]) begin
						controllerinjector_roundrobin7_grant <= 1'd0;
					end else begin
						if (controllerinjector_roundrobin7_request[1]) begin
							controllerinjector_roundrobin7_grant <= 1'd1;
						end else begin
							if (controllerinjector_roundrobin7_request[2]) begin
								controllerinjector_roundrobin7_grant <= 2'd2;
							end else begin
								if (controllerinjector_roundrobin7_request[3]) begin
									controllerinjector_roundrobin7_grant <= 2'd3;
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (controllerinjector_roundrobin7_request[0]) begin
					controllerinjector_roundrobin7_grant <= 1'd0;
				end else begin
					if (controllerinjector_roundrobin7_request[1]) begin
						controllerinjector_roundrobin7_grant <= 1'd1;
					end else begin
						if (controllerinjector_roundrobin7_request[2]) begin
							controllerinjector_roundrobin7_grant <= 2'd2;
						end else begin
							if (controllerinjector_roundrobin7_request[3]) begin
								controllerinjector_roundrobin7_grant <= 2'd3;
							end else begin
								if (controllerinjector_roundrobin7_request[4]) begin
									controllerinjector_roundrobin7_grant <= 3'd4;
								end
							end
						end
					end
				end
			end
		endcase
	end
	hdmi2usbsoc_adr_offset_r <= hdmi2usbsoc_interface0_wb_sdram_adr[0];
	cache_state <= cache_next_state;
	litedramwishbonebridge_state <= litedramwishbonebridge_next_state;
	hdmi2usbsoc_hdmi_in0_edid_sda_drv_reg <= hdmi2usbsoc_hdmi_in0_edid_sda_drv;
	{hdmi2usbsoc_hdmi_in0_edid_samp_carry, hdmi2usbsoc_hdmi_in0_edid_samp_count} <= (hdmi2usbsoc_hdmi_in0_edid_samp_count + 1'd1);
	if (hdmi2usbsoc_hdmi_in0_edid_samp_carry) begin
		hdmi2usbsoc_hdmi_in0_edid_scl_i <= hdmi2usbsoc_hdmi_in0_edid_scl_raw;
		hdmi2usbsoc_hdmi_in0_edid_sda_i <= hdmi2usbsoc_hdmi_in0_edid_sda_raw;
	end
	hdmi2usbsoc_hdmi_in0_edid_scl_r <= hdmi2usbsoc_hdmi_in0_edid_scl_i;
	hdmi2usbsoc_hdmi_in0_edid_sda_r <= hdmi2usbsoc_hdmi_in0_edid_sda_i;
	if (hdmi2usbsoc_hdmi_in0_edid_start) begin
		hdmi2usbsoc_hdmi_in0_edid_counter <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_in0_edid_scl_rising) begin
		if ((hdmi2usbsoc_hdmi_in0_edid_counter == 4'd8)) begin
			hdmi2usbsoc_hdmi_in0_edid_counter <= 1'd0;
		end else begin
			hdmi2usbsoc_hdmi_in0_edid_counter <= (hdmi2usbsoc_hdmi_in0_edid_counter + 1'd1);
			hdmi2usbsoc_hdmi_in0_edid_din <= {hdmi2usbsoc_hdmi_in0_edid_din[6:0], hdmi2usbsoc_hdmi_in0_edid_sda_i};
		end
	end
	if (hdmi2usbsoc_hdmi_in0_edid_update_is_read) begin
		hdmi2usbsoc_hdmi_in0_edid_is_read <= hdmi2usbsoc_hdmi_in0_edid_din[0];
	end
	if (hdmi2usbsoc_hdmi_in0_edid_oc_load) begin
		hdmi2usbsoc_hdmi_in0_edid_offset_counter <= hdmi2usbsoc_hdmi_in0_edid_din;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_edid_oc_inc) begin
			hdmi2usbsoc_hdmi_in0_edid_offset_counter <= (hdmi2usbsoc_hdmi_in0_edid_offset_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in0_edid_data_drv_en) begin
		hdmi2usbsoc_hdmi_in0_edid_data_drv <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_edid_data_drv_stop) begin
			hdmi2usbsoc_hdmi_in0_edid_data_drv <= 1'd0;
		end
	end
	if (hdmi2usbsoc_hdmi_in0_edid_data_drv_en) begin
		case (hdmi2usbsoc_hdmi_in0_edid_counter)
			1'd0: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[7];
			end
			1'd1: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[6];
			end
			2'd2: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[5];
			end
			2'd3: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[4];
			end
			3'd4: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[3];
			end
			3'd5: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[2];
			end
			3'd6: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[1];
			end
			default: begin
				hdmi2usbsoc_hdmi_in0_edid_data_bit <= hdmi2usbsoc_hdmi_in0_edid_dat_r[0];
			end
		endcase
	end
	edid0_state <= edid0_next_state;
	if ((hdmi2usbsoc_hdmi_in0_pll_read_re | hdmi2usbsoc_hdmi_in0_pll_write_re)) begin
		hdmi2usbsoc_hdmi_in0_pll_drdy_status <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_pll_drdy) begin
			hdmi2usbsoc_hdmi_in0_pll_drdy_status <= 1'd1;
		end
	end
	if (((hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_i | hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_i) | hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_master_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_o) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_master_pending <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_i | hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_i) | hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_slave_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_o) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_master_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_slave_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_inc_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_do_delay_dec_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture0_do_reset_lateness_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_wer0_o) begin
		hdmi2usbsoc_hdmi_in0_wer0_wer_counter_sys <= hdmi2usbsoc_hdmi_in0_wer0_wer_counter_r;
	end
	if (hdmi2usbsoc_hdmi_in0_wer0_update_re) begin
		hdmi2usbsoc_hdmi_in0_wer0_status <= hdmi2usbsoc_hdmi_in0_wer0_wer_counter_sys;
	end
	hdmi2usbsoc_hdmi_in0_wer0_toggle_o_r <= hdmi2usbsoc_hdmi_in0_wer0_toggle_o;
	if (((hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_i | hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_i) | hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_master_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_o) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_master_pending <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_i | hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_i) | hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_slave_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_o) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_master_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_slave_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_inc_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_do_delay_dec_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture1_do_reset_lateness_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_wer1_o) begin
		hdmi2usbsoc_hdmi_in0_wer1_wer_counter_sys <= hdmi2usbsoc_hdmi_in0_wer1_wer_counter_r;
	end
	if (hdmi2usbsoc_hdmi_in0_wer1_update_re) begin
		hdmi2usbsoc_hdmi_in0_wer1_status <= hdmi2usbsoc_hdmi_in0_wer1_wer_counter_sys;
	end
	hdmi2usbsoc_hdmi_in0_wer1_toggle_o_r <= hdmi2usbsoc_hdmi_in0_wer1_toggle_o;
	if (((hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_i | hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_i) | hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_master_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_o) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_master_pending <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_i | hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_i) | hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_slave_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_o) begin
			hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_o;
	hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_o_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_master_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_slave_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_inc_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_do_delay_dec_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_i) begin
		hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_i <= (~hdmi2usbsoc_hdmi_in0_s6datacapture2_do_reset_lateness_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in0_wer2_o) begin
		hdmi2usbsoc_hdmi_in0_wer2_wer_counter_sys <= hdmi2usbsoc_hdmi_in0_wer2_wer_counter_r;
	end
	if (hdmi2usbsoc_hdmi_in0_wer2_update_re) begin
		hdmi2usbsoc_hdmi_in0_wer2_status <= hdmi2usbsoc_hdmi_in0_wer2_wer_counter_sys;
	end
	hdmi2usbsoc_hdmi_in0_wer2_toggle_o_r <= hdmi2usbsoc_hdmi_in0_wer2_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_frame_overflow_re) begin
		hdmi2usbsoc_hdmi_in0_frame_overflow_mask <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_o) begin
			hdmi2usbsoc_hdmi_in0_frame_overflow_mask <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_binary <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next_binary;
	hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_next;
	if (hdmi2usbsoc_hdmi_in0_frame_overflow_reset_i) begin
		hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_i <= (~hdmi2usbsoc_hdmi_in0_frame_overflow_reset_toggle_i);
	end
	hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_o_r <= hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_o;
	if (hdmi2usbsoc_hdmi_in0_dma_reset_words) begin
		hdmi2usbsoc_hdmi_in0_dma_current_address <= hdmi2usbsoc_hdmi_in0_dma_slot_array_address;
		hdmi2usbsoc_hdmi_in0_dma_mwords_remaining <= hdmi2usbsoc_hdmi_in0_dma_frame_size_storage;
	end else begin
		if (hdmi2usbsoc_hdmi_in0_dma_count_word) begin
			hdmi2usbsoc_hdmi_in0_dma_current_address <= (hdmi2usbsoc_hdmi_in0_dma_current_address + 1'd1);
			hdmi2usbsoc_hdmi_in0_dma_mwords_remaining <= (hdmi2usbsoc_hdmi_in0_dma_mwords_remaining - 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in0_dma_slot_array_change_slot) begin
		if (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_valid) begin
			hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot <= 1'd1;
		end
		if (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_valid) begin
			hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_we & hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_in0_dma_fifo_replace))) begin
		hdmi2usbsoc_hdmi_in0_dma_fifo_produce <= (hdmi2usbsoc_hdmi_in0_dma_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_in0_dma_fifo_do_read) begin
		hdmi2usbsoc_hdmi_in0_dma_fifo_consume <= (hdmi2usbsoc_hdmi_in0_dma_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_we & hdmi2usbsoc_hdmi_in0_dma_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_in0_dma_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_in0_dma_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_in0_dma_fifo_level <= (hdmi2usbsoc_hdmi_in0_dma_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_in0_dma_fifo_do_read) begin
			hdmi2usbsoc_hdmi_in0_dma_fifo_level <= (hdmi2usbsoc_hdmi_in0_dma_fifo_level - 1'd1);
		end
	end
	dma0_state <= dma0_next_state;
	hdmi2usbsoc_hdmi_in1_edid_sda_drv_reg <= hdmi2usbsoc_hdmi_in1_edid_sda_drv;
	{hdmi2usbsoc_hdmi_in1_edid_samp_carry, hdmi2usbsoc_hdmi_in1_edid_samp_count} <= (hdmi2usbsoc_hdmi_in1_edid_samp_count + 1'd1);
	if (hdmi2usbsoc_hdmi_in1_edid_samp_carry) begin
		hdmi2usbsoc_hdmi_in1_edid_scl_i <= hdmi2usbsoc_hdmi_in1_edid_scl_raw;
		hdmi2usbsoc_hdmi_in1_edid_sda_i <= hdmi2usbsoc_hdmi_in1_edid_sda_raw;
	end
	hdmi2usbsoc_hdmi_in1_edid_scl_r <= hdmi2usbsoc_hdmi_in1_edid_scl_i;
	hdmi2usbsoc_hdmi_in1_edid_sda_r <= hdmi2usbsoc_hdmi_in1_edid_sda_i;
	if (hdmi2usbsoc_hdmi_in1_edid_start) begin
		hdmi2usbsoc_hdmi_in1_edid_counter <= 1'd0;
	end
	if (hdmi2usbsoc_hdmi_in1_edid_scl_rising) begin
		if ((hdmi2usbsoc_hdmi_in1_edid_counter == 4'd8)) begin
			hdmi2usbsoc_hdmi_in1_edid_counter <= 1'd0;
		end else begin
			hdmi2usbsoc_hdmi_in1_edid_counter <= (hdmi2usbsoc_hdmi_in1_edid_counter + 1'd1);
			hdmi2usbsoc_hdmi_in1_edid_din <= {hdmi2usbsoc_hdmi_in1_edid_din[6:0], hdmi2usbsoc_hdmi_in1_edid_sda_i};
		end
	end
	if (hdmi2usbsoc_hdmi_in1_edid_update_is_read) begin
		hdmi2usbsoc_hdmi_in1_edid_is_read <= hdmi2usbsoc_hdmi_in1_edid_din[0];
	end
	if (hdmi2usbsoc_hdmi_in1_edid_oc_load) begin
		hdmi2usbsoc_hdmi_in1_edid_offset_counter <= hdmi2usbsoc_hdmi_in1_edid_din;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_edid_oc_inc) begin
			hdmi2usbsoc_hdmi_in1_edid_offset_counter <= (hdmi2usbsoc_hdmi_in1_edid_offset_counter + 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in1_edid_data_drv_en) begin
		hdmi2usbsoc_hdmi_in1_edid_data_drv <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_edid_data_drv_stop) begin
			hdmi2usbsoc_hdmi_in1_edid_data_drv <= 1'd0;
		end
	end
	if (hdmi2usbsoc_hdmi_in1_edid_data_drv_en) begin
		case (hdmi2usbsoc_hdmi_in1_edid_counter)
			1'd0: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[7];
			end
			1'd1: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[6];
			end
			2'd2: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[5];
			end
			2'd3: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[4];
			end
			3'd4: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[3];
			end
			3'd5: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[2];
			end
			3'd6: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[1];
			end
			default: begin
				hdmi2usbsoc_hdmi_in1_edid_data_bit <= hdmi2usbsoc_hdmi_in1_edid_dat_r[0];
			end
		endcase
	end
	edid1_state <= edid1_next_state;
	if ((hdmi2usbsoc_hdmi_in1_pll_read_re | hdmi2usbsoc_hdmi_in1_pll_write_re)) begin
		hdmi2usbsoc_hdmi_in1_pll_drdy_status <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_pll_drdy) begin
			hdmi2usbsoc_hdmi_in1_pll_drdy_status <= 1'd1;
		end
	end
	if (((hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_i | hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_i) | hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_master_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_o) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_master_pending <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_i | hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_i) | hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_slave_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_o) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_master_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_slave_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_inc_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_do_delay_dec_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture0_do_reset_lateness_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_wer0_o) begin
		hdmi2usbsoc_hdmi_in1_wer0_wer_counter_sys <= hdmi2usbsoc_hdmi_in1_wer0_wer_counter_r;
	end
	if (hdmi2usbsoc_hdmi_in1_wer0_update_re) begin
		hdmi2usbsoc_hdmi_in1_wer0_status <= hdmi2usbsoc_hdmi_in1_wer0_wer_counter_sys;
	end
	hdmi2usbsoc_hdmi_in1_wer0_toggle_o_r <= hdmi2usbsoc_hdmi_in1_wer0_toggle_o;
	if (((hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_i | hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_i) | hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_master_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_o) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_master_pending <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_i | hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_i) | hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_slave_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_o) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_master_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_slave_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_inc_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_do_delay_dec_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture1_do_reset_lateness_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_wer1_o) begin
		hdmi2usbsoc_hdmi_in1_wer1_wer_counter_sys <= hdmi2usbsoc_hdmi_in1_wer1_wer_counter_r;
	end
	if (hdmi2usbsoc_hdmi_in1_wer1_update_re) begin
		hdmi2usbsoc_hdmi_in1_wer1_status <= hdmi2usbsoc_hdmi_in1_wer1_wer_counter_sys;
	end
	hdmi2usbsoc_hdmi_in1_wer1_toggle_o_r <= hdmi2usbsoc_hdmi_in1_wer1_toggle_o;
	if (((hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_i | hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_i) | hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_master_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_o) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_master_pending <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_i | hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_i) | hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_i)) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_slave_pending <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_o) begin
			hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_slave_pending <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_o;
	hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_o_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_master_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_cal_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_slave_rst_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_inc_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_do_delay_dec_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_i) begin
		hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_i <= (~hdmi2usbsoc_hdmi_in1_s6datacapture2_do_reset_lateness_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_in1_wer2_o) begin
		hdmi2usbsoc_hdmi_in1_wer2_wer_counter_sys <= hdmi2usbsoc_hdmi_in1_wer2_wer_counter_r;
	end
	if (hdmi2usbsoc_hdmi_in1_wer2_update_re) begin
		hdmi2usbsoc_hdmi_in1_wer2_status <= hdmi2usbsoc_hdmi_in1_wer2_wer_counter_sys;
	end
	hdmi2usbsoc_hdmi_in1_wer2_toggle_o_r <= hdmi2usbsoc_hdmi_in1_wer2_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_frame_overflow_re) begin
		hdmi2usbsoc_hdmi_in1_frame_overflow_mask <= 1'd1;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_o) begin
			hdmi2usbsoc_hdmi_in1_frame_overflow_mask <= 1'd0;
		end
	end
	hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_binary <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next_binary;
	hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_next;
	if (hdmi2usbsoc_hdmi_in1_frame_overflow_reset_i) begin
		hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_i <= (~hdmi2usbsoc_hdmi_in1_frame_overflow_reset_toggle_i);
	end
	hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_o_r <= hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_o;
	if (hdmi2usbsoc_hdmi_in1_dma_reset_words) begin
		hdmi2usbsoc_hdmi_in1_dma_current_address <= hdmi2usbsoc_hdmi_in1_dma_slot_array_address;
		hdmi2usbsoc_hdmi_in1_dma_mwords_remaining <= hdmi2usbsoc_hdmi_in1_dma_frame_size_storage;
	end else begin
		if (hdmi2usbsoc_hdmi_in1_dma_count_word) begin
			hdmi2usbsoc_hdmi_in1_dma_current_address <= (hdmi2usbsoc_hdmi_in1_dma_current_address + 1'd1);
			hdmi2usbsoc_hdmi_in1_dma_mwords_remaining <= (hdmi2usbsoc_hdmi_in1_dma_mwords_remaining - 1'd1);
		end
	end
	if (hdmi2usbsoc_hdmi_in1_dma_slot_array_change_slot) begin
		if (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_valid) begin
			hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot <= 1'd1;
		end
		if (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_valid) begin
			hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot <= 1'd0;
		end
	end
	if (((hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_we & hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_in1_dma_fifo_replace))) begin
		hdmi2usbsoc_hdmi_in1_dma_fifo_produce <= (hdmi2usbsoc_hdmi_in1_dma_fifo_produce + 1'd1);
	end
	if (hdmi2usbsoc_hdmi_in1_dma_fifo_do_read) begin
		hdmi2usbsoc_hdmi_in1_dma_fifo_consume <= (hdmi2usbsoc_hdmi_in1_dma_fifo_consume + 1'd1);
	end
	if (((hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_we & hdmi2usbsoc_hdmi_in1_dma_fifo_syncfifo_writable) & (~hdmi2usbsoc_hdmi_in1_dma_fifo_replace))) begin
		if ((~hdmi2usbsoc_hdmi_in1_dma_fifo_do_read)) begin
			hdmi2usbsoc_hdmi_in1_dma_fifo_level <= (hdmi2usbsoc_hdmi_in1_dma_fifo_level + 1'd1);
		end
	end else begin
		if (hdmi2usbsoc_hdmi_in1_dma_fifo_do_read) begin
			hdmi2usbsoc_hdmi_in1_dma_fifo_level <= (hdmi2usbsoc_hdmi_in1_dma_fifo_level - 1'd1);
		end
	end
	dma1_state <= dma1_next_state;
	hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary;
	hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_next;
	if (hdmi2usbsoc_hdmi_out0_core_i) begin
		hdmi2usbsoc_hdmi_out0_core_toggle_i <= (~hdmi2usbsoc_hdmi_out0_core_toggle_i);
	end
	if (hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_remaining_bits <= 4'd10;
		hdmi2usbsoc_hdmi_out0_driver_clocking_sr <= hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage;
	end else begin
		if (hdmi2usbsoc_hdmi_out0_driver_clocking_transmitting) begin
			hdmi2usbsoc_hdmi_out0_driver_clocking_remaining_bits <= (hdmi2usbsoc_hdmi_out0_driver_clocking_remaining_bits - 1'd1);
			hdmi2usbsoc_hdmi_out0_driver_clocking_sr <= hdmi2usbsoc_hdmi_out0_driver_clocking_sr[9:1];
		end
	end
	if (hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_busy_counter <= 4'd13;
	end else begin
		if (hdmi2usbsoc_hdmi_out0_driver_clocking_busy) begin
			hdmi2usbsoc_hdmi_out0_driver_clocking_busy_counter <= (hdmi2usbsoc_hdmi_out0_driver_clocking_busy_counter - 1'd1);
		end
	end
	if ((hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_re | hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_re)) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy_status <= 1'd0;
	end else begin
		if (hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy) begin
			hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy_status <= 1'd1;
		end
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_binary <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next_binary;
	hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_next;
	if (hdmi2usbsoc_hdmi_out1_core_i) begin
		hdmi2usbsoc_hdmi_out1_core_toggle_i <= (~hdmi2usbsoc_hdmi_out1_core_toggle_i);
	end
	if ((encoder_reader_start_r & encoder_reader_start_re)) begin
		encoder_reader_base <= encoder_reader_base_storage;
	end
	if (encoder_reader_h_clr) begin
		encoder_reader_h <= 1'd0;
	end else begin
		if (encoder_reader_h_clr_lsb) begin
			encoder_reader_h[2:0] <= 1'd0;
			encoder_reader_h[15:3] <= encoder_reader_h[15:3];
		end else begin
			if (encoder_reader_h_inc) begin
				encoder_reader_h <= encoder_reader_h_next;
			end
		end
	end
	if (encoder_reader_v_clr) begin
		encoder_reader_v <= 1'd0;
	end else begin
		if (encoder_reader_v_inc) begin
			encoder_reader_v <= (encoder_reader_v + 1'd1);
		end else begin
			if (encoder_reader_v_dec7) begin
				encoder_reader_v <= (encoder_reader_v - 3'd7);
			end
		end
	end
	if (encoder_reader_request_issued) begin
		if ((~encoder_reader_data_dequeued)) begin
			encoder_reader_rsv_level <= (encoder_reader_rsv_level + 1'd1);
		end
	end else begin
		if (encoder_reader_data_dequeued) begin
			encoder_reader_rsv_level <= (encoder_reader_rsv_level - 1'd1);
		end
	end
	if (((encoder_reader_fifo_syncfifo_we & encoder_reader_fifo_syncfifo_writable) & (~encoder_reader_fifo_replace))) begin
		encoder_reader_fifo_produce <= (encoder_reader_fifo_produce + 1'd1);
	end
	if (encoder_reader_fifo_do_read) begin
		encoder_reader_fifo_consume <= (encoder_reader_fifo_consume + 1'd1);
	end
	if (((encoder_reader_fifo_syncfifo_we & encoder_reader_fifo_syncfifo_writable) & (~encoder_reader_fifo_replace))) begin
		if ((~encoder_reader_fifo_do_read)) begin
			encoder_reader_fifo_level <= (encoder_reader_fifo_level + 1'd1);
		end
	end else begin
		if (encoder_reader_fifo_do_read) begin
			encoder_reader_fifo_level <= (encoder_reader_fifo_level - 1'd1);
		end
	end
	encoderdmareader_state <= encoderdmareader_next_state;
	encoder_cdc_graycounter0_q_binary <= encoder_cdc_graycounter0_q_next_binary;
	encoder_cdc_graycounter0_q <= encoder_cdc_graycounter0_q_next;
	case (hdmi2usbsoc_grant)
		1'd0: begin
			if ((~hdmi2usbsoc_request[0])) begin
				if (hdmi2usbsoc_request[1]) begin
					hdmi2usbsoc_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~hdmi2usbsoc_request[1])) begin
				if (hdmi2usbsoc_request[0]) begin
					hdmi2usbsoc_grant <= 1'd0;
				end
			end
		end
	endcase
	hdmi2usbsoc_slave_sel_r <= hdmi2usbsoc_slave_sel;
	hdmi2usbsoc_interface0_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank0_sel) begin
		case (hdmi2usbsoc_interface0_bank_bus_adr[3:0])
			1'd0: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_base3_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_base2_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_base1_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_base0_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_h_width1_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_h_width0_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_v_width1_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_v_width0_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= encoder_reader_start_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface0_bank_bus_dat_r <= hdmi2usbsoc_csrbank0_done_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank0_base3_re) begin
		encoder_reader_base_storage_full[31:24] <= hdmi2usbsoc_csrbank0_base3_r;
	end
	if (hdmi2usbsoc_csrbank0_base2_re) begin
		encoder_reader_base_storage_full[23:16] <= hdmi2usbsoc_csrbank0_base2_r;
	end
	if (hdmi2usbsoc_csrbank0_base1_re) begin
		encoder_reader_base_storage_full[15:8] <= hdmi2usbsoc_csrbank0_base1_r;
	end
	if (hdmi2usbsoc_csrbank0_base0_re) begin
		encoder_reader_base_storage_full[7:0] <= hdmi2usbsoc_csrbank0_base0_r;
	end
	encoder_reader_base_re <= hdmi2usbsoc_csrbank0_base0_re;
	if (hdmi2usbsoc_csrbank0_h_width1_re) begin
		encoder_reader_h_width_storage_full[15:8] <= hdmi2usbsoc_csrbank0_h_width1_r;
	end
	if (hdmi2usbsoc_csrbank0_h_width0_re) begin
		encoder_reader_h_width_storage_full[7:0] <= hdmi2usbsoc_csrbank0_h_width0_r;
	end
	encoder_reader_h_width_re <= hdmi2usbsoc_csrbank0_h_width0_re;
	if (hdmi2usbsoc_csrbank0_v_width1_re) begin
		encoder_reader_v_width_storage_full[15:8] <= hdmi2usbsoc_csrbank0_v_width1_r;
	end
	if (hdmi2usbsoc_csrbank0_v_width0_re) begin
		encoder_reader_v_width_storage_full[7:0] <= hdmi2usbsoc_csrbank0_v_width0_r;
	end
	encoder_reader_v_width_re <= hdmi2usbsoc_csrbank0_v_width0_re;
	hdmi2usbsoc_sram0_sel_r <= hdmi2usbsoc_sram0_sel;
	hdmi2usbsoc_interface1_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank1_sel) begin
		case (hdmi2usbsoc_interface1_bank_bus_adr[6:0])
			1'd0: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_edid_hpd_notif_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_edid_hpd_en0_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_pll_reset0_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_locked_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_pll_adr0_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_pll_dat_r1_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_pll_dat_r0_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_pll_read_w;
			end
			4'd10: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_pll_write_w;
			end
			4'd11: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_clocking_pll_drdy_w;
			end
			4'd12: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_dly_ctl_w;
			end
			4'd13: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data0_cap_dly_busy_w;
			end
			4'd14: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data0_cap_phase_w;
			end
			4'd15: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_s6datacapture0_phase_reset_w;
			end
			5'd16: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data0_charsync_char_synced_w;
			end
			5'd17: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data0_charsync_ctl_pos_w;
			end
			5'd18: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_wer0_update_w;
			end
			5'd19: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data0_wer_value2_w;
			end
			5'd20: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data0_wer_value1_w;
			end
			5'd21: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data0_wer_value0_w;
			end
			5'd22: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_dly_ctl_w;
			end
			5'd23: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data1_cap_dly_busy_w;
			end
			5'd24: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data1_cap_phase_w;
			end
			5'd25: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_s6datacapture1_phase_reset_w;
			end
			5'd26: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data1_charsync_char_synced_w;
			end
			5'd27: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data1_charsync_ctl_pos_w;
			end
			5'd28: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_wer1_update_w;
			end
			5'd29: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data1_wer_value2_w;
			end
			5'd30: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data1_wer_value1_w;
			end
			5'd31: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data1_wer_value0_w;
			end
			6'd32: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_dly_ctl_w;
			end
			6'd33: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data2_cap_dly_busy_w;
			end
			6'd34: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data2_cap_phase_w;
			end
			6'd35: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_s6datacapture2_phase_reset_w;
			end
			6'd36: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data2_charsync_char_synced_w;
			end
			6'd37: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data2_charsync_ctl_pos_w;
			end
			6'd38: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_wer2_update_w;
			end
			6'd39: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data2_wer_value2_w;
			end
			6'd40: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data2_wer_value1_w;
			end
			6'd41: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_data2_wer_value0_w;
			end
			6'd42: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_chansync_channels_synced_w;
			end
			6'd43: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_resdetection_hres1_w;
			end
			6'd44: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_resdetection_hres0_w;
			end
			6'd45: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_resdetection_vres1_w;
			end
			6'd46: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_resdetection_vres0_w;
			end
			6'd47: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_frame_overflow_w;
			end
			6'd48: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_frame_size3_w;
			end
			6'd49: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_frame_size2_w;
			end
			6'd50: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_frame_size1_w;
			end
			6'd51: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_frame_size0_w;
			end
			6'd52: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot0_status0_w;
			end
			6'd53: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot0_address3_w;
			end
			6'd54: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot0_address2_w;
			end
			6'd55: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot0_address1_w;
			end
			6'd56: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot0_address0_w;
			end
			6'd57: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot1_status0_w;
			end
			6'd58: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot1_address3_w;
			end
			6'd59: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot1_address2_w;
			end
			6'd60: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot1_address1_w;
			end
			6'd61: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_slot1_address0_w;
			end
			6'd62: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_dma_slot_array_status_w;
			end
			6'd63: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in0_dma_slot_array_pending_w;
			end
			7'd64: begin
				hdmi2usbsoc_interface1_bank_bus_dat_r <= hdmi2usbsoc_csrbank1_dma_ev_enable0_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank1_edid_hpd_en0_re) begin
		hdmi2usbsoc_hdmi_in0_edid_storage_full <= hdmi2usbsoc_csrbank1_edid_hpd_en0_r;
	end
	hdmi2usbsoc_hdmi_in0_edid_re <= hdmi2usbsoc_csrbank1_edid_hpd_en0_re;
	if (hdmi2usbsoc_csrbank1_clocking_pll_reset0_re) begin
		hdmi2usbsoc_hdmi_in0_pll_reset_storage_full <= hdmi2usbsoc_csrbank1_clocking_pll_reset0_r;
	end
	hdmi2usbsoc_hdmi_in0_pll_reset_re <= hdmi2usbsoc_csrbank1_clocking_pll_reset0_re;
	if (hdmi2usbsoc_csrbank1_clocking_pll_adr0_re) begin
		hdmi2usbsoc_hdmi_in0_pll_adr_storage_full[4:0] <= hdmi2usbsoc_csrbank1_clocking_pll_adr0_r;
	end
	hdmi2usbsoc_hdmi_in0_pll_adr_re <= hdmi2usbsoc_csrbank1_clocking_pll_adr0_re;
	if (hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_re) begin
		hdmi2usbsoc_hdmi_in0_pll_dat_w_storage_full[15:8] <= hdmi2usbsoc_csrbank1_clocking_pll_dat_w1_r;
	end
	if (hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_re) begin
		hdmi2usbsoc_hdmi_in0_pll_dat_w_storage_full[7:0] <= hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_r;
	end
	hdmi2usbsoc_hdmi_in0_pll_dat_w_re <= hdmi2usbsoc_csrbank1_clocking_pll_dat_w0_re;
	if (hdmi2usbsoc_csrbank1_dma_frame_size3_re) begin
		hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[26:24] <= hdmi2usbsoc_csrbank1_dma_frame_size3_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_frame_size2_re) begin
		hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[23:16] <= hdmi2usbsoc_csrbank1_dma_frame_size2_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_frame_size1_re) begin
		hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[15:8] <= hdmi2usbsoc_csrbank1_dma_frame_size1_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_frame_size0_re) begin
		hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full[7:0] <= hdmi2usbsoc_csrbank1_dma_frame_size0_r;
	end
	hdmi2usbsoc_hdmi_in0_dma_frame_size_re <= hdmi2usbsoc_csrbank1_dma_frame_size0_re;
	if (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_we) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage_full <= (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_dat_w <<< 1'd0);
	end
	if (hdmi2usbsoc_csrbank1_dma_slot0_status0_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage_full[1:0] <= hdmi2usbsoc_csrbank1_dma_slot0_status0_r;
	end
	hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_re <= hdmi2usbsoc_csrbank1_dma_slot0_status0_re;
	if (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_we) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full <= (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_dat_w <<< 2'd3);
	end
	if (hdmi2usbsoc_csrbank1_dma_slot0_address3_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[26:24] <= hdmi2usbsoc_csrbank1_dma_slot0_address3_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_slot0_address2_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[23:16] <= hdmi2usbsoc_csrbank1_dma_slot0_address2_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_slot0_address1_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[15:8] <= hdmi2usbsoc_csrbank1_dma_slot0_address1_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_slot0_address0_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full[7:0] <= hdmi2usbsoc_csrbank1_dma_slot0_address0_r;
	end
	hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_re <= hdmi2usbsoc_csrbank1_dma_slot0_address0_re;
	if (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_we) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage_full <= (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_dat_w <<< 1'd0);
	end
	if (hdmi2usbsoc_csrbank1_dma_slot1_status0_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage_full[1:0] <= hdmi2usbsoc_csrbank1_dma_slot1_status0_r;
	end
	hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_re <= hdmi2usbsoc_csrbank1_dma_slot1_status0_re;
	if (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_we) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full <= (hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_dat_w <<< 2'd3);
	end
	if (hdmi2usbsoc_csrbank1_dma_slot1_address3_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[26:24] <= hdmi2usbsoc_csrbank1_dma_slot1_address3_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_slot1_address2_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[23:16] <= hdmi2usbsoc_csrbank1_dma_slot1_address2_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_slot1_address1_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[15:8] <= hdmi2usbsoc_csrbank1_dma_slot1_address1_r;
	end
	if (hdmi2usbsoc_csrbank1_dma_slot1_address0_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full[7:0] <= hdmi2usbsoc_csrbank1_dma_slot1_address0_r;
	end
	hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_re <= hdmi2usbsoc_csrbank1_dma_slot1_address0_re;
	if (hdmi2usbsoc_csrbank1_dma_ev_enable0_re) begin
		hdmi2usbsoc_hdmi_in0_dma_slot_array_storage_full[1:0] <= hdmi2usbsoc_csrbank1_dma_ev_enable0_r;
	end
	hdmi2usbsoc_hdmi_in0_dma_slot_array_re <= hdmi2usbsoc_csrbank1_dma_ev_enable0_re;
	hdmi2usbsoc_sram1_sel_r <= hdmi2usbsoc_sram1_sel;
	hdmi2usbsoc_interface2_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank2_sel) begin
		case (hdmi2usbsoc_interface2_bank_bus_adr[6:0])
			1'd0: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_edid_hpd_notif_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_edid_hpd_en0_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_pll_reset0_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_locked_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_pll_adr0_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_pll_dat_r1_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_pll_dat_r0_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_pll_read_w;
			end
			4'd10: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_pll_write_w;
			end
			4'd11: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_clocking_pll_drdy_w;
			end
			4'd12: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_dly_ctl_w;
			end
			4'd13: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data0_cap_dly_busy_w;
			end
			4'd14: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data0_cap_phase_w;
			end
			4'd15: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_s6datacapture0_phase_reset_w;
			end
			5'd16: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data0_charsync_char_synced_w;
			end
			5'd17: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data0_charsync_ctl_pos_w;
			end
			5'd18: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_wer0_update_w;
			end
			5'd19: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data0_wer_value2_w;
			end
			5'd20: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data0_wer_value1_w;
			end
			5'd21: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data0_wer_value0_w;
			end
			5'd22: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_dly_ctl_w;
			end
			5'd23: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data1_cap_dly_busy_w;
			end
			5'd24: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data1_cap_phase_w;
			end
			5'd25: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_s6datacapture1_phase_reset_w;
			end
			5'd26: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data1_charsync_char_synced_w;
			end
			5'd27: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data1_charsync_ctl_pos_w;
			end
			5'd28: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_wer1_update_w;
			end
			5'd29: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data1_wer_value2_w;
			end
			5'd30: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data1_wer_value1_w;
			end
			5'd31: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data1_wer_value0_w;
			end
			6'd32: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_dly_ctl_w;
			end
			6'd33: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data2_cap_dly_busy_w;
			end
			6'd34: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data2_cap_phase_w;
			end
			6'd35: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_s6datacapture2_phase_reset_w;
			end
			6'd36: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data2_charsync_char_synced_w;
			end
			6'd37: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data2_charsync_ctl_pos_w;
			end
			6'd38: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_wer2_update_w;
			end
			6'd39: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data2_wer_value2_w;
			end
			6'd40: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data2_wer_value1_w;
			end
			6'd41: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_data2_wer_value0_w;
			end
			6'd42: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_chansync_channels_synced_w;
			end
			6'd43: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_resdetection_hres1_w;
			end
			6'd44: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_resdetection_hres0_w;
			end
			6'd45: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_resdetection_vres1_w;
			end
			6'd46: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_resdetection_vres0_w;
			end
			6'd47: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_frame_overflow_w;
			end
			6'd48: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_frame_size3_w;
			end
			6'd49: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_frame_size2_w;
			end
			6'd50: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_frame_size1_w;
			end
			6'd51: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_frame_size0_w;
			end
			6'd52: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot0_status0_w;
			end
			6'd53: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot0_address3_w;
			end
			6'd54: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot0_address2_w;
			end
			6'd55: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot0_address1_w;
			end
			6'd56: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot0_address0_w;
			end
			6'd57: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot1_status0_w;
			end
			6'd58: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot1_address3_w;
			end
			6'd59: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot1_address2_w;
			end
			6'd60: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot1_address1_w;
			end
			6'd61: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_slot1_address0_w;
			end
			6'd62: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_dma_slot_array_status_w;
			end
			6'd63: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_hdmi_in1_dma_slot_array_pending_w;
			end
			7'd64: begin
				hdmi2usbsoc_interface2_bank_bus_dat_r <= hdmi2usbsoc_csrbank2_dma_ev_enable0_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank2_edid_hpd_en0_re) begin
		hdmi2usbsoc_hdmi_in1_edid_storage_full <= hdmi2usbsoc_csrbank2_edid_hpd_en0_r;
	end
	hdmi2usbsoc_hdmi_in1_edid_re <= hdmi2usbsoc_csrbank2_edid_hpd_en0_re;
	if (hdmi2usbsoc_csrbank2_clocking_pll_reset0_re) begin
		hdmi2usbsoc_hdmi_in1_pll_reset_storage_full <= hdmi2usbsoc_csrbank2_clocking_pll_reset0_r;
	end
	hdmi2usbsoc_hdmi_in1_pll_reset_re <= hdmi2usbsoc_csrbank2_clocking_pll_reset0_re;
	if (hdmi2usbsoc_csrbank2_clocking_pll_adr0_re) begin
		hdmi2usbsoc_hdmi_in1_pll_adr_storage_full[4:0] <= hdmi2usbsoc_csrbank2_clocking_pll_adr0_r;
	end
	hdmi2usbsoc_hdmi_in1_pll_adr_re <= hdmi2usbsoc_csrbank2_clocking_pll_adr0_re;
	if (hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_re) begin
		hdmi2usbsoc_hdmi_in1_pll_dat_w_storage_full[15:8] <= hdmi2usbsoc_csrbank2_clocking_pll_dat_w1_r;
	end
	if (hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_re) begin
		hdmi2usbsoc_hdmi_in1_pll_dat_w_storage_full[7:0] <= hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_r;
	end
	hdmi2usbsoc_hdmi_in1_pll_dat_w_re <= hdmi2usbsoc_csrbank2_clocking_pll_dat_w0_re;
	if (hdmi2usbsoc_csrbank2_dma_frame_size3_re) begin
		hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[26:24] <= hdmi2usbsoc_csrbank2_dma_frame_size3_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_frame_size2_re) begin
		hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[23:16] <= hdmi2usbsoc_csrbank2_dma_frame_size2_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_frame_size1_re) begin
		hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[15:8] <= hdmi2usbsoc_csrbank2_dma_frame_size1_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_frame_size0_re) begin
		hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full[7:0] <= hdmi2usbsoc_csrbank2_dma_frame_size0_r;
	end
	hdmi2usbsoc_hdmi_in1_dma_frame_size_re <= hdmi2usbsoc_csrbank2_dma_frame_size0_re;
	if (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_we) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage_full <= (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_dat_w <<< 1'd0);
	end
	if (hdmi2usbsoc_csrbank2_dma_slot0_status0_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage_full[1:0] <= hdmi2usbsoc_csrbank2_dma_slot0_status0_r;
	end
	hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_re <= hdmi2usbsoc_csrbank2_dma_slot0_status0_re;
	if (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_we) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full <= (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_dat_w <<< 2'd3);
	end
	if (hdmi2usbsoc_csrbank2_dma_slot0_address3_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[26:24] <= hdmi2usbsoc_csrbank2_dma_slot0_address3_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_slot0_address2_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[23:16] <= hdmi2usbsoc_csrbank2_dma_slot0_address2_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_slot0_address1_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[15:8] <= hdmi2usbsoc_csrbank2_dma_slot0_address1_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_slot0_address0_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full[7:0] <= hdmi2usbsoc_csrbank2_dma_slot0_address0_r;
	end
	hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_re <= hdmi2usbsoc_csrbank2_dma_slot0_address0_re;
	if (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_we) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage_full <= (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_dat_w <<< 1'd0);
	end
	if (hdmi2usbsoc_csrbank2_dma_slot1_status0_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage_full[1:0] <= hdmi2usbsoc_csrbank2_dma_slot1_status0_r;
	end
	hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_re <= hdmi2usbsoc_csrbank2_dma_slot1_status0_re;
	if (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_we) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full <= (hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_dat_w <<< 2'd3);
	end
	if (hdmi2usbsoc_csrbank2_dma_slot1_address3_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[26:24] <= hdmi2usbsoc_csrbank2_dma_slot1_address3_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_slot1_address2_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[23:16] <= hdmi2usbsoc_csrbank2_dma_slot1_address2_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_slot1_address1_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[15:8] <= hdmi2usbsoc_csrbank2_dma_slot1_address1_r;
	end
	if (hdmi2usbsoc_csrbank2_dma_slot1_address0_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full[7:0] <= hdmi2usbsoc_csrbank2_dma_slot1_address0_r;
	end
	hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_re <= hdmi2usbsoc_csrbank2_dma_slot1_address0_re;
	if (hdmi2usbsoc_csrbank2_dma_ev_enable0_re) begin
		hdmi2usbsoc_hdmi_in1_dma_slot_array_storage_full[1:0] <= hdmi2usbsoc_csrbank2_dma_ev_enable0_r;
	end
	hdmi2usbsoc_hdmi_in1_dma_slot_array_re <= hdmi2usbsoc_csrbank2_dma_ev_enable0_re;
	hdmi2usbsoc_interface3_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank3_sel) begin
		case (hdmi2usbsoc_interface3_bank_bus_adr[5:0])
			1'd0: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_underflow_enable0_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_hdmi_out0_core_underflow_update_underflow_update_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_underflow_counter3_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_underflow_counter2_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_underflow_counter1_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_underflow_counter0_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_enable0_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hres1_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hres0_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_w;
			end
			4'd10: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_w;
			end
			4'd11: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_w;
			end
			4'd12: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_w;
			end
			4'd13: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hscan1_w;
			end
			4'd14: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_hscan0_w;
			end
			4'd15: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vres1_w;
			end
			5'd16: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vres0_w;
			end
			5'd17: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_w;
			end
			5'd18: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_w;
			end
			5'd19: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_w;
			end
			5'd20: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_w;
			end
			5'd21: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vscan1_w;
			end
			5'd22: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_vscan0_w;
			end
			5'd23: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_base3_w;
			end
			5'd24: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_base2_w;
			end
			5'd25: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_base1_w;
			end
			5'd26: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_base0_w;
			end
			5'd27: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_length3_w;
			end
			5'd28: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_length2_w;
			end
			5'd29: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_length1_w;
			end
			5'd30: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_core_initiator_length0_w;
			end
			5'd31: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_w;
			end
			6'd32: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_w;
			end
			6'd33: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_hdmi_out0_driver_clocking_send_cmd_data_w;
			end
			6'd34: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_hdmi_out0_driver_clocking_send_go_w;
			end
			6'd35: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_status_w;
			end
			6'd36: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_w;
			end
			6'd37: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_w;
			end
			6'd38: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r1_w;
			end
			6'd39: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_r0_w;
			end
			6'd40: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_w;
			end
			6'd41: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_w;
			end
			6'd42: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_w;
			end
			6'd43: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_w;
			end
			6'd44: begin
				hdmi2usbsoc_interface3_bank_bus_dat_r <= hdmi2usbsoc_csrbank3_driver_clocking_pll_drdy_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank3_core_underflow_enable0_re) begin
		hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage_full <= hdmi2usbsoc_csrbank3_core_underflow_enable0_r;
	end
	hdmi2usbsoc_hdmi_out0_core_underflow_enable_re <= hdmi2usbsoc_csrbank3_core_underflow_enable0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_enable0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage_full <= hdmi2usbsoc_csrbank3_core_initiator_enable0_r;
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_enable_re <= hdmi2usbsoc_csrbank3_core_initiator_enable0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_hres1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_hres_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_hres1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_hres0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_hres_backstore, hdmi2usbsoc_csrbank3_core_initiator_hres0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_re <= hdmi2usbsoc_csrbank3_core_initiator_hres0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_hsync_start_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_hsync_start1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_hsync_start_backstore, hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_re <= hdmi2usbsoc_csrbank3_core_initiator_hsync_start0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_hsync_end_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_hsync_end1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_hsync_end_backstore, hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_re <= hdmi2usbsoc_csrbank3_core_initiator_hsync_end0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_hscan1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_hscan_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_hscan1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_hscan0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_hscan_backstore, hdmi2usbsoc_csrbank3_core_initiator_hscan0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_re <= hdmi2usbsoc_csrbank3_core_initiator_hscan0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_vres1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_vres_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_vres1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_vres0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_vres_backstore, hdmi2usbsoc_csrbank3_core_initiator_vres0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_re <= hdmi2usbsoc_csrbank3_core_initiator_vres0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_vsync_start_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_vsync_start1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_vsync_start_backstore, hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_re <= hdmi2usbsoc_csrbank3_core_initiator_vsync_start0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_vsync_end_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_vsync_end1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_vsync_end_backstore, hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_re <= hdmi2usbsoc_csrbank3_core_initiator_vsync_end0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_vscan1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_vscan_backstore[3:0] <= hdmi2usbsoc_csrbank3_core_initiator_vscan1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_vscan0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_vscan_backstore, hdmi2usbsoc_csrbank3_core_initiator_vscan0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_re <= hdmi2usbsoc_csrbank3_core_initiator_vscan0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_base3_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_base_backstore[23:16] <= hdmi2usbsoc_csrbank3_core_initiator_base3_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_base2_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_base_backstore[15:8] <= hdmi2usbsoc_csrbank3_core_initiator_base2_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_base1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_base_backstore[7:0] <= hdmi2usbsoc_csrbank3_core_initiator_base1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_base0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_base_backstore, hdmi2usbsoc_csrbank3_core_initiator_base0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_re <= hdmi2usbsoc_csrbank3_core_initiator_base0_re;
	if (hdmi2usbsoc_csrbank3_core_initiator_length3_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_length_backstore[23:16] <= hdmi2usbsoc_csrbank3_core_initiator_length3_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_length2_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_length_backstore[15:8] <= hdmi2usbsoc_csrbank3_core_initiator_length2_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_length1_re) begin
		hdmi2usbsoc_csrbank3_core_initiator_length_backstore[7:0] <= hdmi2usbsoc_csrbank3_core_initiator_length1_r;
	end
	if (hdmi2usbsoc_csrbank3_core_initiator_length0_re) begin
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full <= {hdmi2usbsoc_csrbank3_core_initiator_length_backstore, hdmi2usbsoc_csrbank3_core_initiator_length0_r};
	end
	hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_re <= hdmi2usbsoc_csrbank3_core_initiator_length0_re;
	if (hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage_full[9:8] <= hdmi2usbsoc_csrbank3_driver_clocking_cmd_data1_r;
	end
	if (hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage_full[7:0] <= hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_r;
	end
	hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_re <= hdmi2usbsoc_csrbank3_driver_clocking_cmd_data0_re;
	if (hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage_full <= hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_r;
	end
	hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_re <= hdmi2usbsoc_csrbank3_driver_clocking_pll_reset0_re;
	if (hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage_full[4:0] <= hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_r;
	end
	hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_re <= hdmi2usbsoc_csrbank3_driver_clocking_pll_adr0_re;
	if (hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage_full[15:8] <= hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w1_r;
	end
	if (hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_re) begin
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage_full[7:0] <= hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_r;
	end
	hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_re <= hdmi2usbsoc_csrbank3_driver_clocking_pll_dat_w0_re;
	hdmi2usbsoc_interface4_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank4_sel) begin
		case (hdmi2usbsoc_interface4_bank_bus_adr[4:0])
			1'd0: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_underflow_enable0_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_hdmi_out1_core_underflow_update_underflow_update_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_underflow_counter3_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_underflow_counter2_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_underflow_counter1_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_underflow_counter0_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_enable0_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hres1_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hres0_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_w;
			end
			4'd10: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_w;
			end
			4'd11: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_w;
			end
			4'd12: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_w;
			end
			4'd13: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hscan1_w;
			end
			4'd14: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_hscan0_w;
			end
			4'd15: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vres1_w;
			end
			5'd16: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vres0_w;
			end
			5'd17: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_w;
			end
			5'd18: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_w;
			end
			5'd19: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_w;
			end
			5'd20: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_w;
			end
			5'd21: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vscan1_w;
			end
			5'd22: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_vscan0_w;
			end
			5'd23: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_base3_w;
			end
			5'd24: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_base2_w;
			end
			5'd25: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_base1_w;
			end
			5'd26: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_base0_w;
			end
			5'd27: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_length3_w;
			end
			5'd28: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_length2_w;
			end
			5'd29: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_length1_w;
			end
			5'd30: begin
				hdmi2usbsoc_interface4_bank_bus_dat_r <= hdmi2usbsoc_csrbank4_core_initiator_length0_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank4_core_underflow_enable0_re) begin
		hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage_full <= hdmi2usbsoc_csrbank4_core_underflow_enable0_r;
	end
	hdmi2usbsoc_hdmi_out1_core_underflow_enable_re <= hdmi2usbsoc_csrbank4_core_underflow_enable0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_enable0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage_full <= hdmi2usbsoc_csrbank4_core_initiator_enable0_r;
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_enable_re <= hdmi2usbsoc_csrbank4_core_initiator_enable0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_hres1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_hres_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_hres1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_hres0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_hres_backstore, hdmi2usbsoc_csrbank4_core_initiator_hres0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_re <= hdmi2usbsoc_csrbank4_core_initiator_hres0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_hsync_start_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_hsync_start1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_hsync_start_backstore, hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_re <= hdmi2usbsoc_csrbank4_core_initiator_hsync_start0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_hsync_end_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_hsync_end1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_hsync_end_backstore, hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_re <= hdmi2usbsoc_csrbank4_core_initiator_hsync_end0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_hscan1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_hscan_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_hscan1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_hscan0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_hscan_backstore, hdmi2usbsoc_csrbank4_core_initiator_hscan0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_re <= hdmi2usbsoc_csrbank4_core_initiator_hscan0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_vres1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_vres_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_vres1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_vres0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_vres_backstore, hdmi2usbsoc_csrbank4_core_initiator_vres0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_re <= hdmi2usbsoc_csrbank4_core_initiator_vres0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_vsync_start_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_vsync_start1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_vsync_start_backstore, hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_re <= hdmi2usbsoc_csrbank4_core_initiator_vsync_start0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_vsync_end_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_vsync_end1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_vsync_end_backstore, hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_re <= hdmi2usbsoc_csrbank4_core_initiator_vsync_end0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_vscan1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_vscan_backstore[3:0] <= hdmi2usbsoc_csrbank4_core_initiator_vscan1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_vscan0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_vscan_backstore, hdmi2usbsoc_csrbank4_core_initiator_vscan0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_re <= hdmi2usbsoc_csrbank4_core_initiator_vscan0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_base3_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_base_backstore[23:16] <= hdmi2usbsoc_csrbank4_core_initiator_base3_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_base2_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_base_backstore[15:8] <= hdmi2usbsoc_csrbank4_core_initiator_base2_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_base1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_base_backstore[7:0] <= hdmi2usbsoc_csrbank4_core_initiator_base1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_base0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_base_backstore, hdmi2usbsoc_csrbank4_core_initiator_base0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_re <= hdmi2usbsoc_csrbank4_core_initiator_base0_re;
	if (hdmi2usbsoc_csrbank4_core_initiator_length3_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_length_backstore[23:16] <= hdmi2usbsoc_csrbank4_core_initiator_length3_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_length2_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_length_backstore[15:8] <= hdmi2usbsoc_csrbank4_core_initiator_length2_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_length1_re) begin
		hdmi2usbsoc_csrbank4_core_initiator_length_backstore[7:0] <= hdmi2usbsoc_csrbank4_core_initiator_length1_r;
	end
	if (hdmi2usbsoc_csrbank4_core_initiator_length0_re) begin
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full <= {hdmi2usbsoc_csrbank4_core_initiator_length_backstore, hdmi2usbsoc_csrbank4_core_initiator_length0_r};
	end
	hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_re <= hdmi2usbsoc_csrbank4_core_initiator_length0_re;
	hdmi2usbsoc_sram2_sel_r <= hdmi2usbsoc_sram2_sel;
	hdmi2usbsoc_interface5_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank5_sel) begin
		case (hdmi2usbsoc_interface5_bank_bus_adr[5:0])
			1'd0: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id7_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id6_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id5_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id4_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id3_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id2_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id1_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_dna_id0_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit19_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit18_w;
			end
			4'd10: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit17_w;
			end
			4'd11: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit16_w;
			end
			4'd12: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit15_w;
			end
			4'd13: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit14_w;
			end
			4'd14: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit13_w;
			end
			4'd15: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit12_w;
			end
			5'd16: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit11_w;
			end
			5'd17: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit10_w;
			end
			5'd18: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit9_w;
			end
			5'd19: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit8_w;
			end
			5'd20: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit7_w;
			end
			5'd21: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit6_w;
			end
			5'd22: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit5_w;
			end
			5'd23: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit4_w;
			end
			5'd24: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit3_w;
			end
			5'd25: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit2_w;
			end
			5'd26: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit1_w;
			end
			5'd27: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_git_commit0_w;
			end
			5'd28: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform7_w;
			end
			5'd29: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform6_w;
			end
			5'd30: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform5_w;
			end
			5'd31: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform4_w;
			end
			6'd32: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform3_w;
			end
			6'd33: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform2_w;
			end
			6'd34: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform1_w;
			end
			6'd35: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_platform0_w;
			end
			6'd36: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target7_w;
			end
			6'd37: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target6_w;
			end
			6'd38: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target5_w;
			end
			6'd39: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target4_w;
			end
			6'd40: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target3_w;
			end
			6'd41: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target2_w;
			end
			6'd42: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target1_w;
			end
			6'd43: begin
				hdmi2usbsoc_interface5_bank_bus_dat_r <= hdmi2usbsoc_csrbank5_platform_target0_w;
			end
		endcase
	end
	hdmi2usbsoc_interface6_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank6_sel) begin
		case (hdmi2usbsoc_interface6_bank_bus_adr[5:0])
			1'd0: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_control0_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_command0_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_sdram_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_address1_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_address0_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_w;
			end
			4'd10: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_rddata3_w;
			end
			4'd11: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_rddata2_w;
			end
			4'd12: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_rddata1_w;
			end
			4'd13: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi0_rddata0_w;
			end
			4'd14: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_command0_w;
			end
			4'd15: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_sdram_phaseinjector1_command_issue_w;
			end
			5'd16: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_address1_w;
			end
			5'd17: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_address0_w;
			end
			5'd18: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_w;
			end
			5'd19: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_w;
			end
			5'd20: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_w;
			end
			5'd21: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_w;
			end
			5'd22: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_w;
			end
			5'd23: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_rddata3_w;
			end
			5'd24: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_rddata2_w;
			end
			5'd25: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_rddata1_w;
			end
			5'd26: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_dfii_pi1_rddata0_w;
			end
			5'd27: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_sdram_bandwidth_update_w;
			end
			5'd28: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_controller_bandwidth_nreads2_w;
			end
			5'd29: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_controller_bandwidth_nreads1_w;
			end
			5'd30: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_controller_bandwidth_nreads0_w;
			end
			5'd31: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites2_w;
			end
			6'd32: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites1_w;
			end
			6'd33: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_controller_bandwidth_nwrites0_w;
			end
			6'd34: begin
				hdmi2usbsoc_interface6_bank_bus_dat_r <= hdmi2usbsoc_csrbank6_controller_bandwidth_data_width_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank6_dfii_control0_re) begin
		hdmi2usbsoc_sdram_storage_full[3:0] <= hdmi2usbsoc_csrbank6_dfii_control0_r;
	end
	hdmi2usbsoc_sdram_re <= hdmi2usbsoc_csrbank6_dfii_control0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi0_command0_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_command_storage_full[5:0] <= hdmi2usbsoc_csrbank6_dfii_pi0_command0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector0_command_re <= hdmi2usbsoc_csrbank6_dfii_pi0_command0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi0_address1_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_address_storage_full[12:8] <= hdmi2usbsoc_csrbank6_dfii_pi0_address1_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi0_address0_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_address_storage_full[7:0] <= hdmi2usbsoc_csrbank6_dfii_pi0_address0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector0_address_re <= hdmi2usbsoc_csrbank6_dfii_pi0_address0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_baddress_storage_full[2:0] <= hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector0_baddress_re <= hdmi2usbsoc_csrbank6_dfii_pi0_baddress0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[31:24] <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata3_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[23:16] <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata2_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[15:8] <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata1_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_re) begin
		hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full[7:0] <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector0_wrdata_re <= hdmi2usbsoc_csrbank6_dfii_pi0_wrdata0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi1_command0_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_command_storage_full[5:0] <= hdmi2usbsoc_csrbank6_dfii_pi1_command0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector1_command_re <= hdmi2usbsoc_csrbank6_dfii_pi1_command0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi1_address1_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_address_storage_full[12:8] <= hdmi2usbsoc_csrbank6_dfii_pi1_address1_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi1_address0_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_address_storage_full[7:0] <= hdmi2usbsoc_csrbank6_dfii_pi1_address0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector1_address_re <= hdmi2usbsoc_csrbank6_dfii_pi1_address0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_baddress_storage_full[2:0] <= hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector1_baddress_re <= hdmi2usbsoc_csrbank6_dfii_pi1_baddress0_re;
	if (hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[31:24] <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata3_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[23:16] <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata2_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[15:8] <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata1_r;
	end
	if (hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_re) begin
		hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full[7:0] <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_r;
	end
	hdmi2usbsoc_sdram_phaseinjector1_wrdata_re <= hdmi2usbsoc_csrbank6_dfii_pi1_wrdata0_re;
	hdmi2usbsoc_interface7_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank7_sel) begin
		case (hdmi2usbsoc_interface7_bank_bus_adr[1:0])
			1'd0: begin
				hdmi2usbsoc_interface7_bank_bus_dat_r <= hdmi2usbsoc_csrbank7_bitbang0_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface7_bank_bus_dat_r <= hdmi2usbsoc_csrbank7_miso_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface7_bank_bus_dat_r <= hdmi2usbsoc_csrbank7_bitbang_en0_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank7_bitbang0_re) begin
		hdmi2usbsoc_bitbang_storage_full[3:0] <= hdmi2usbsoc_csrbank7_bitbang0_r;
	end
	hdmi2usbsoc_bitbang_re <= hdmi2usbsoc_csrbank7_bitbang0_re;
	if (hdmi2usbsoc_csrbank7_bitbang_en0_re) begin
		hdmi2usbsoc_bitbang_en_storage_full <= hdmi2usbsoc_csrbank7_bitbang_en0_r;
	end
	hdmi2usbsoc_bitbang_en_re <= hdmi2usbsoc_csrbank7_bitbang_en0_re;
	hdmi2usbsoc_interface8_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank8_sel) begin
		case (hdmi2usbsoc_interface8_bank_bus_adr[4:0])
			1'd0: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_load3_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_load2_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_load1_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_load0_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_reload3_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_reload2_w;
			end
			3'd6: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_reload1_w;
			end
			3'd7: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_reload0_w;
			end
			4'd8: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_en0_w;
			end
			4'd9: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_hdmi2usbsoc_timer0_update_value_w;
			end
			4'd10: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_value3_w;
			end
			4'd11: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_value2_w;
			end
			4'd12: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_value1_w;
			end
			4'd13: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_value0_w;
			end
			4'd14: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_status_w;
			end
			4'd15: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_pending_w;
			end
			5'd16: begin
				hdmi2usbsoc_interface8_bank_bus_dat_r <= hdmi2usbsoc_csrbank8_ev_enable0_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank8_load3_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[31:24] <= hdmi2usbsoc_csrbank8_load3_r;
	end
	if (hdmi2usbsoc_csrbank8_load2_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[23:16] <= hdmi2usbsoc_csrbank8_load2_r;
	end
	if (hdmi2usbsoc_csrbank8_load1_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[15:8] <= hdmi2usbsoc_csrbank8_load1_r;
	end
	if (hdmi2usbsoc_csrbank8_load0_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full[7:0] <= hdmi2usbsoc_csrbank8_load0_r;
	end
	hdmi2usbsoc_hdmi2usbsoc_timer0_load_re <= hdmi2usbsoc_csrbank8_load0_re;
	if (hdmi2usbsoc_csrbank8_reload3_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[31:24] <= hdmi2usbsoc_csrbank8_reload3_r;
	end
	if (hdmi2usbsoc_csrbank8_reload2_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[23:16] <= hdmi2usbsoc_csrbank8_reload2_r;
	end
	if (hdmi2usbsoc_csrbank8_reload1_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[15:8] <= hdmi2usbsoc_csrbank8_reload1_r;
	end
	if (hdmi2usbsoc_csrbank8_reload0_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full[7:0] <= hdmi2usbsoc_csrbank8_reload0_r;
	end
	hdmi2usbsoc_hdmi2usbsoc_timer0_reload_re <= hdmi2usbsoc_csrbank8_reload0_re;
	if (hdmi2usbsoc_csrbank8_en0_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage_full <= hdmi2usbsoc_csrbank8_en0_r;
	end
	hdmi2usbsoc_hdmi2usbsoc_timer0_en_re <= hdmi2usbsoc_csrbank8_en0_re;
	if (hdmi2usbsoc_csrbank8_ev_enable0_re) begin
		hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage_full <= hdmi2usbsoc_csrbank8_ev_enable0_r;
	end
	hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_re <= hdmi2usbsoc_csrbank8_ev_enable0_re;
	hdmi2usbsoc_interface9_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank9_sel) begin
		case (hdmi2usbsoc_interface9_bank_bus_adr[2:0])
			1'd0: begin
				hdmi2usbsoc_interface9_bank_bus_dat_r <= hdmi2usbsoc_hdmi2usbsoc_uart_rxtx_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface9_bank_bus_dat_r <= hdmi2usbsoc_csrbank9_txfull_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface9_bank_bus_dat_r <= hdmi2usbsoc_csrbank9_rxempty_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface9_bank_bus_dat_r <= hdmi2usbsoc_hdmi2usbsoc_uart_status_w;
			end
			3'd4: begin
				hdmi2usbsoc_interface9_bank_bus_dat_r <= hdmi2usbsoc_hdmi2usbsoc_uart_pending_w;
			end
			3'd5: begin
				hdmi2usbsoc_interface9_bank_bus_dat_r <= hdmi2usbsoc_csrbank9_ev_enable0_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank9_ev_enable0_re) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_storage_full[1:0] <= hdmi2usbsoc_csrbank9_ev_enable0_r;
	end
	hdmi2usbsoc_hdmi2usbsoc_uart_re <= hdmi2usbsoc_csrbank9_ev_enable0_re;
	hdmi2usbsoc_interface10_bank_bus_dat_r <= 1'd0;
	if (hdmi2usbsoc_csrbank10_sel) begin
		case (hdmi2usbsoc_interface10_bank_bus_adr[1:0])
			1'd0: begin
				hdmi2usbsoc_interface10_bank_bus_dat_r <= hdmi2usbsoc_csrbank10_tuning_word3_w;
			end
			1'd1: begin
				hdmi2usbsoc_interface10_bank_bus_dat_r <= hdmi2usbsoc_csrbank10_tuning_word2_w;
			end
			2'd2: begin
				hdmi2usbsoc_interface10_bank_bus_dat_r <= hdmi2usbsoc_csrbank10_tuning_word1_w;
			end
			2'd3: begin
				hdmi2usbsoc_interface10_bank_bus_dat_r <= hdmi2usbsoc_csrbank10_tuning_word0_w;
			end
		endcase
	end
	if (hdmi2usbsoc_csrbank10_tuning_word3_re) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[31:24] <= hdmi2usbsoc_csrbank10_tuning_word3_r;
	end
	if (hdmi2usbsoc_csrbank10_tuning_word2_re) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[23:16] <= hdmi2usbsoc_csrbank10_tuning_word2_r;
	end
	if (hdmi2usbsoc_csrbank10_tuning_word1_re) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[15:8] <= hdmi2usbsoc_csrbank10_tuning_word1_r;
	end
	if (hdmi2usbsoc_csrbank10_tuning_word0_re) begin
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full[7:0] <= hdmi2usbsoc_csrbank10_tuning_word0_r;
	end
	hdmi2usbsoc_hdmi2usbsoc_uart_phy_re <= hdmi2usbsoc_csrbank10_tuning_word0_re;
	if (sys_rst) begin
		hdmi2usbsoc_hdmi2usbsoc_rom_bus_ack <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_sram_bus_ack <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_interface_adr <= 14'd0;
		hdmi2usbsoc_hdmi2usbsoc_interface_we <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_interface_dat_w <= 8'd0;
		hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_dat_r <= 32'd0;
		hdmi2usbsoc_hdmi2usbsoc_bus_wishbone_ack <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_counter <= 2'd0;
		serial_tx <= 1'd1;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_storage_full <= 32'd6597069;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_re <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_sink_ready <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_txen <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_tx <= 32'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_reg <= 8'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_bitcount <= 4'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_tx_busy <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_valid <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_source_payload_data <= 8'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_uart_clk_rxen <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_phase_accumulator_rx <= 32'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_r <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_reg <= 8'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_bitcount <= 4'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_phy_rx_busy <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_pending <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_old_trigger <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_pending <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_old_trigger <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_storage_full <= 2'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_re <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_level <= 5'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_produce <= 4'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_consume <= 4'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_level <= 5'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_produce <= 4'd0;
		hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_consume <= 4'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_load_storage_full <= 32'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_load_re <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_reload_storage_full <= 32'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_reload_re <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_en_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_en_re <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_value_status <= 32'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_zero_pending <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_zero_old_trigger <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_eventmanager_re <= 1'd0;
		hdmi2usbsoc_hdmi2usbsoc_timer0_value <= 32'd0;
		hdmi2usbsoc_dna_status <= 57'd0;
		hdmi2usbsoc_dna_cnt <= 7'd0;
		hdmi2usbsoc_bus_ack <= 1'd0;
		hdmi2usbsoc_bitbang_storage_full <= 4'd0;
		hdmi2usbsoc_bitbang_re <= 1'd0;
		hdmi2usbsoc_bitbang_en_storage_full <= 1'd0;
		hdmi2usbsoc_bitbang_en_re <= 1'd0;
		hdmi2usbsoc_cs_n <= 1'd1;
		hdmi2usbsoc_clk <= 1'd0;
		hdmi2usbsoc_dq_oe <= 1'd0;
		hdmi2usbsoc_sr <= 32'd0;
		hdmi2usbsoc_i1 <= 2'd0;
		hdmi2usbsoc_dqi <= 4'd0;
		hdmi2usbsoc_counter <= 8'd0;
		hdmi2usbsoc_ddrphy_phase_sys <= 1'd0;
		hdmi2usbsoc_ddrphy_bitslip_cnt <= 4'd0;
		hdmi2usbsoc_ddrphy_bitslip_inc <= 1'd0;
		hdmi2usbsoc_ddrphy_record2_wrdata <= 32'd0;
		hdmi2usbsoc_ddrphy_record2_wrdata_mask <= 4'd0;
		hdmi2usbsoc_ddrphy_record3_wrdata <= 32'd0;
		hdmi2usbsoc_ddrphy_record3_wrdata_mask <= 4'd0;
		hdmi2usbsoc_ddrphy_drive_dq_n1 <= 1'd0;
		hdmi2usbsoc_ddrphy_wrdata_en_d <= 1'd0;
		hdmi2usbsoc_ddrphy_rddata_sr <= 5'd0;
		hdmi2usbsoc_sdram_storage_full <= 4'd0;
		hdmi2usbsoc_sdram_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector0_command_storage_full <= 6'd0;
		hdmi2usbsoc_sdram_phaseinjector0_command_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector0_address_storage_full <= 13'd0;
		hdmi2usbsoc_sdram_phaseinjector0_address_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector0_baddress_storage_full <= 3'd0;
		hdmi2usbsoc_sdram_phaseinjector0_baddress_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector0_wrdata_storage_full <= 32'd0;
		hdmi2usbsoc_sdram_phaseinjector0_wrdata_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector0_status <= 32'd0;
		hdmi2usbsoc_sdram_phaseinjector1_command_storage_full <= 6'd0;
		hdmi2usbsoc_sdram_phaseinjector1_command_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector1_address_storage_full <= 13'd0;
		hdmi2usbsoc_sdram_phaseinjector1_address_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector1_baddress_storage_full <= 3'd0;
		hdmi2usbsoc_sdram_phaseinjector1_baddress_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector1_wrdata_storage_full <= 32'd0;
		hdmi2usbsoc_sdram_phaseinjector1_wrdata_re <= 1'd0;
		hdmi2usbsoc_sdram_phaseinjector1_status <= 32'd0;
		hdmi2usbsoc_sdram_dfi_p0_address <= 13'd0;
		hdmi2usbsoc_sdram_dfi_p0_bank <= 3'd0;
		hdmi2usbsoc_sdram_dfi_p0_cas_n <= 1'd1;
		hdmi2usbsoc_sdram_dfi_p0_ras_n <= 1'd1;
		hdmi2usbsoc_sdram_dfi_p0_we_n <= 1'd1;
		hdmi2usbsoc_sdram_dfi_p0_wrdata_en <= 1'd0;
		hdmi2usbsoc_sdram_dfi_p0_rddata_en <= 1'd0;
		hdmi2usbsoc_sdram_dfi_p1_address <= 13'd0;
		hdmi2usbsoc_sdram_dfi_p1_bank <= 3'd0;
		hdmi2usbsoc_sdram_dfi_p1_cas_n <= 1'd1;
		hdmi2usbsoc_sdram_dfi_p1_ras_n <= 1'd1;
		hdmi2usbsoc_sdram_dfi_p1_we_n <= 1'd1;
		hdmi2usbsoc_sdram_dfi_p1_wrdata_en <= 1'd0;
		hdmi2usbsoc_sdram_dfi_p1_rddata_en <= 1'd0;
		hdmi2usbsoc_sdram_cmd_payload_a <= 13'd0;
		hdmi2usbsoc_sdram_cmd_payload_ba <= 3'd0;
		hdmi2usbsoc_sdram_cmd_payload_cas <= 1'd0;
		hdmi2usbsoc_sdram_cmd_payload_ras <= 1'd0;
		hdmi2usbsoc_sdram_cmd_payload_we <= 1'd0;
		hdmi2usbsoc_sdram_seq_done <= 1'd0;
		hdmi2usbsoc_sdram_counter <= 4'd0;
		hdmi2usbsoc_sdram_count <= 10'd585;
		hdmi2usbsoc_sdram_bankmachine0_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine0_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine0_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine0_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine0_count <= 3'd4;
		hdmi2usbsoc_sdram_bankmachine1_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine1_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine1_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine1_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine1_count <= 3'd4;
		hdmi2usbsoc_sdram_bankmachine2_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine2_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine2_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine2_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine2_count <= 3'd4;
		hdmi2usbsoc_sdram_bankmachine3_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine3_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine3_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine3_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine3_count <= 3'd4;
		hdmi2usbsoc_sdram_bankmachine4_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine4_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine4_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine4_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine4_count <= 3'd4;
		hdmi2usbsoc_sdram_bankmachine5_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine5_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine5_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine5_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine5_count <= 3'd4;
		hdmi2usbsoc_sdram_bankmachine6_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine6_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine6_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine6_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine6_count <= 3'd4;
		hdmi2usbsoc_sdram_bankmachine7_level <= 4'd0;
		hdmi2usbsoc_sdram_bankmachine7_produce <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine7_consume <= 3'd0;
		hdmi2usbsoc_sdram_bankmachine7_has_openrow <= 1'd0;
		hdmi2usbsoc_sdram_bankmachine7_count <= 3'd4;
		hdmi2usbsoc_sdram_choose_cmd_grant <= 3'd0;
		hdmi2usbsoc_sdram_choose_req_grant <= 3'd0;
		hdmi2usbsoc_sdram_time0 <= 5'd0;
		hdmi2usbsoc_sdram_time1 <= 4'd0;
		hdmi2usbsoc_sdram_bandwidth_nreads_status <= 24'd0;
		hdmi2usbsoc_sdram_bandwidth_nwrites_status <= 24'd0;
		hdmi2usbsoc_sdram_bandwidth_cmd_valid <= 1'd0;
		hdmi2usbsoc_sdram_bandwidth_cmd_ready <= 1'd0;
		hdmi2usbsoc_sdram_bandwidth_cmd_is_read <= 1'd0;
		hdmi2usbsoc_sdram_bandwidth_cmd_is_write <= 1'd0;
		hdmi2usbsoc_sdram_bandwidth_counter <= 24'd0;
		hdmi2usbsoc_sdram_bandwidth_period <= 1'd0;
		hdmi2usbsoc_sdram_bandwidth_nreads <= 24'd0;
		hdmi2usbsoc_sdram_bandwidth_nwrites <= 24'd0;
		hdmi2usbsoc_sdram_bandwidth_nreads_r <= 24'd0;
		hdmi2usbsoc_sdram_bandwidth_nwrites_r <= 24'd0;
		hdmi2usbsoc_adr_offset_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_sda_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_sda_drv_reg <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_scl_i <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_samp_count <= 6'd0;
		hdmi2usbsoc_hdmi_in0_edid_samp_carry <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_scl_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_sda_r <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_din <= 8'd0;
		hdmi2usbsoc_hdmi_in0_edid_counter <= 4'd0;
		hdmi2usbsoc_hdmi_in0_edid_is_read <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_offset_counter <= 7'd0;
		hdmi2usbsoc_hdmi_in0_edid_data_bit <= 1'd0;
		hdmi2usbsoc_hdmi_in0_edid_data_drv <= 1'd0;
		hdmi2usbsoc_hdmi_in0_pll_reset_storage_full <= 1'd1;
		hdmi2usbsoc_hdmi_in0_pll_reset_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_pll_adr_storage_full <= 5'd0;
		hdmi2usbsoc_hdmi_in0_pll_adr_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_pll_dat_w_storage_full <= 16'd0;
		hdmi2usbsoc_hdmi_in0_pll_dat_w_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_pll_drdy_status <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture0_sys_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer0_status <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer0_wer_counter_sys <= 24'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture1_sys_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer1_status <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer1_wer_counter_sys <= 24'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_s6datacapture2_sys_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in0_wer2_status <= 24'd0;
		hdmi2usbsoc_hdmi_in0_wer2_wer_counter_sys <= 24'd0;
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q <= 10'd0;
		hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter1_q_binary <= 10'd0;
		hdmi2usbsoc_hdmi_in0_frame_overflow_mask <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_frame_size_storage_full <= 27'd0;
		hdmi2usbsoc_hdmi_in0_dma_frame_size_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_storage_full <= 2'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_status_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_storage_full <= 27'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot0_address_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_storage_full <= 2'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_status_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_storage_full <= 27'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_slot1_address_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_storage_full <= 2'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_re <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_slot_array_current_slot <= 1'd0;
		hdmi2usbsoc_hdmi_in0_dma_current_address <= 24'd0;
		hdmi2usbsoc_hdmi_in0_dma_mwords_remaining <= 24'd0;
		hdmi2usbsoc_hdmi_in0_dma_fifo_level <= 5'd0;
		hdmi2usbsoc_hdmi_in0_dma_fifo_produce <= 4'd0;
		hdmi2usbsoc_hdmi_in0_dma_fifo_consume <= 4'd0;
		hdmi2usbsoc_hdmi_in1_edid_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_sda_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_sda_drv_reg <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_scl_i <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_samp_count <= 6'd0;
		hdmi2usbsoc_hdmi_in1_edid_samp_carry <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_scl_r <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_sda_r <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_din <= 8'd0;
		hdmi2usbsoc_hdmi_in1_edid_counter <= 4'd0;
		hdmi2usbsoc_hdmi_in1_edid_is_read <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_offset_counter <= 7'd0;
		hdmi2usbsoc_hdmi_in1_edid_data_bit <= 1'd0;
		hdmi2usbsoc_hdmi_in1_edid_data_drv <= 1'd0;
		hdmi2usbsoc_hdmi_in1_pll_reset_storage_full <= 1'd1;
		hdmi2usbsoc_hdmi_in1_pll_reset_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_pll_adr_storage_full <= 5'd0;
		hdmi2usbsoc_hdmi_in1_pll_adr_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_pll_dat_w_storage_full <= 16'd0;
		hdmi2usbsoc_hdmi_in1_pll_dat_w_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_pll_drdy_status <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture0_sys_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer0_status <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer0_wer_counter_sys <= 24'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture1_sys_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer1_status <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer1_wer_counter_sys <= 24'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_master_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_s6datacapture2_sys_delay_slave_pending <= 1'd0;
		hdmi2usbsoc_hdmi_in1_wer2_status <= 24'd0;
		hdmi2usbsoc_hdmi_in1_wer2_wer_counter_sys <= 24'd0;
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q <= 10'd0;
		hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter1_q_binary <= 10'd0;
		hdmi2usbsoc_hdmi_in1_frame_overflow_mask <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_frame_size_storage_full <= 27'd0;
		hdmi2usbsoc_hdmi_in1_dma_frame_size_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_storage_full <= 2'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_status_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_storage_full <= 27'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot0_address_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_storage_full <= 2'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_status_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_storage_full <= 27'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_slot1_address_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_storage_full <= 2'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_re <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_slot_array_current_slot <= 1'd0;
		hdmi2usbsoc_hdmi_in1_dma_current_address <= 24'd0;
		hdmi2usbsoc_hdmi_in1_dma_mwords_remaining <= 24'd0;
		hdmi2usbsoc_hdmi_in1_dma_fifo_level <= 5'd0;
		hdmi2usbsoc_hdmi_in1_dma_fifo_produce <= 4'd0;
		hdmi2usbsoc_hdmi_in1_dma_fifo_consume <= 4'd0;
		hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q <= 3'd0;
		hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter1_q_binary <= 3'd0;
		hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q <= 5'd0;
		hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter0_q_binary <= 5'd0;
		hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_underflow_enable_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q <= 2'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary <= 2'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_enable_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_enable_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage0_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage1_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage2_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage3_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage4_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage5_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage6_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage7_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_storage_full <= 32'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage8_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_storage_full <= 32'd0;
		hdmi2usbsoc_hdmi_out0_core_initiator_csrstorage9_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_storage_full <= 10'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_cmd_data_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage_full <= 5'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage_full <= 16'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_re <= 1'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy_status <= 1'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_remaining_bits <= 4'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_sr <= 10'd0;
		hdmi2usbsoc_hdmi_out0_driver_clocking_busy_counter <= 4'd0;
		hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q <= 3'd0;
		hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter3_q_binary <= 3'd0;
		hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q <= 5'd0;
		hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter2_q_binary <= 5'd0;
		hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_underflow_enable_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q <= 2'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter0_q_binary <= 2'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_enable_storage_full <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_enable_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage0_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage1_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage2_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage3_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage4_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage5_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage6_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_storage_full <= 12'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage7_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_storage_full <= 32'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage8_re <= 1'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_storage_full <= 32'd0;
		hdmi2usbsoc_hdmi_out1_core_initiator_csrstorage9_re <= 1'd0;
		encoder_port_counter <= 1'd0;
		encoder_port_converter_source_first <= 1'd0;
		encoder_port_converter_source_last <= 1'd0;
		encoder_port_converter_source_payload_data <= 128'd0;
		encoder_port_converter_source_payload_valid_token_count <= 2'd0;
		encoder_port_converter_demux <= 1'd0;
		encoder_port_converter_strobe_all <= 1'd0;
		encoder_reader_base_storage_full <= 32'd0;
		encoder_reader_base_re <= 1'd0;
		encoder_reader_h_width_storage_full <= 16'd0;
		encoder_reader_h_width_re <= 1'd0;
		encoder_reader_v_width_storage_full <= 16'd0;
		encoder_reader_v_width_re <= 1'd0;
		encoder_reader_rsv_level <= 5'd0;
		encoder_reader_fifo_level <= 5'd0;
		encoder_reader_fifo_produce <= 4'd0;
		encoder_reader_fifo_consume <= 4'd0;
		encoder_reader_base <= 32'd0;
		encoder_reader_h <= 16'd0;
		encoder_reader_v <= 16'd0;
		encoder_cdc_graycounter0_q <= 3'd0;
		encoder_cdc_graycounter0_q_binary <= 3'd0;
		controllerinjector_refresher_state <= 2'd0;
		controllerinjector_bankmachine0_state <= 3'd0;
		controllerinjector_bankmachine1_state <= 3'd0;
		controllerinjector_bankmachine2_state <= 3'd0;
		controllerinjector_bankmachine3_state <= 3'd0;
		controllerinjector_bankmachine4_state <= 3'd0;
		controllerinjector_bankmachine5_state <= 3'd0;
		controllerinjector_bankmachine6_state <= 3'd0;
		controllerinjector_bankmachine7_state <= 3'd0;
		controllerinjector_multiplexer_state <= 4'd0;
		controllerinjector_state <= 1'd0;
		controllerinjector_roundrobin0_grant <= 3'd0;
		controllerinjector_roundrobin1_grant <= 3'd0;
		controllerinjector_roundrobin2_grant <= 3'd0;
		controllerinjector_roundrobin3_grant <= 3'd0;
		controllerinjector_roundrobin4_grant <= 3'd0;
		controllerinjector_roundrobin5_grant <= 3'd0;
		controllerinjector_roundrobin6_grant <= 3'd0;
		controllerinjector_roundrobin7_grant <= 3'd0;
		controllerinjector_new_master_wdata_ready0 <= 1'd0;
		controllerinjector_new_master_wdata_ready1 <= 1'd0;
		controllerinjector_new_master_wdata_ready2 <= 1'd0;
		controllerinjector_new_master_wdata_ready3 <= 1'd0;
		controllerinjector_new_master_wdata_ready4 <= 1'd0;
		controllerinjector_new_master_wdata_ready5 <= 1'd0;
		controllerinjector_new_master_rdata_valid0 <= 1'd0;
		controllerinjector_new_master_rdata_valid1 <= 1'd0;
		controllerinjector_new_master_rdata_valid2 <= 1'd0;
		controllerinjector_new_master_rdata_valid3 <= 1'd0;
		controllerinjector_new_master_rdata_valid4 <= 1'd0;
		controllerinjector_new_master_rdata_valid5 <= 1'd0;
		controllerinjector_new_master_rdata_valid6 <= 1'd0;
		controllerinjector_new_master_rdata_valid7 <= 1'd0;
		controllerinjector_new_master_rdata_valid8 <= 1'd0;
		controllerinjector_new_master_rdata_valid9 <= 1'd0;
		controllerinjector_new_master_rdata_valid10 <= 1'd0;
		controllerinjector_new_master_rdata_valid11 <= 1'd0;
		controllerinjector_new_master_rdata_valid12 <= 1'd0;
		controllerinjector_new_master_rdata_valid13 <= 1'd0;
		controllerinjector_new_master_rdata_valid14 <= 1'd0;
		controllerinjector_new_master_rdata_valid15 <= 1'd0;
		controllerinjector_new_master_rdata_valid16 <= 1'd0;
		controllerinjector_new_master_rdata_valid17 <= 1'd0;
		controllerinjector_new_master_rdata_valid18 <= 1'd0;
		controllerinjector_new_master_rdata_valid19 <= 1'd0;
		controllerinjector_new_master_rdata_valid20 <= 1'd0;
		controllerinjector_new_master_rdata_valid21 <= 1'd0;
		controllerinjector_new_master_rdata_valid22 <= 1'd0;
		controllerinjector_new_master_rdata_valid23 <= 1'd0;
		controllerinjector_new_master_rdata_valid24 <= 1'd0;
		controllerinjector_new_master_rdata_valid25 <= 1'd0;
		controllerinjector_new_master_rdata_valid26 <= 1'd0;
		controllerinjector_new_master_rdata_valid27 <= 1'd0;
		controllerinjector_new_master_rdata_valid28 <= 1'd0;
		controllerinjector_new_master_rdata_valid29 <= 1'd0;
		controllerinjector_new_master_rdata_valid30 <= 1'd0;
		controllerinjector_new_master_rdata_valid31 <= 1'd0;
		controllerinjector_new_master_rdata_valid32 <= 1'd0;
		controllerinjector_new_master_rdata_valid33 <= 1'd0;
		controllerinjector_new_master_rdata_valid34 <= 1'd0;
		controllerinjector_new_master_rdata_valid35 <= 1'd0;
		cache_state <= 3'd0;
		litedramwishbonebridge_state <= 2'd0;
		edid0_state <= 4'd0;
		dma0_state <= 2'd0;
		edid1_state <= 4'd0;
		dma1_state <= 2'd0;
		encoderdmareader_state <= 1'd0;
		hdmi2usbsoc_grant <= 1'd0;
		hdmi2usbsoc_slave_sel_r <= 6'd0;
		hdmi2usbsoc_interface0_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_sram0_sel_r <= 1'd0;
		hdmi2usbsoc_interface1_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_sram1_sel_r <= 1'd0;
		hdmi2usbsoc_interface2_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_interface3_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_csrbank3_core_initiator_hres_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_hsync_start_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_hsync_end_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_hscan_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_vres_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_vsync_start_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_vsync_end_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_vscan_backstore <= 4'd0;
		hdmi2usbsoc_csrbank3_core_initiator_base_backstore <= 24'd0;
		hdmi2usbsoc_csrbank3_core_initiator_length_backstore <= 24'd0;
		hdmi2usbsoc_interface4_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_csrbank4_core_initiator_hres_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_hsync_start_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_hsync_end_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_hscan_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_vres_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_vsync_start_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_vsync_end_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_vscan_backstore <= 4'd0;
		hdmi2usbsoc_csrbank4_core_initiator_base_backstore <= 24'd0;
		hdmi2usbsoc_csrbank4_core_initiator_length_backstore <= 24'd0;
		hdmi2usbsoc_sram2_sel_r <= 1'd0;
		hdmi2usbsoc_interface5_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_interface6_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_interface7_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_interface8_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_interface9_bank_bus_dat_r <= 8'd0;
		hdmi2usbsoc_interface10_bank_bus_dat_r <= 8'd0;
	end
	xilinxmultiregimpl0_regs0 <= serial_rx;
	xilinxmultiregimpl0_regs1 <= xilinxmultiregimpl0_regs0;
	xilinxmultiregimpl1_regs0 <= hdmi_in0_scl;
	xilinxmultiregimpl1_regs1 <= xilinxmultiregimpl1_regs0;
	xilinxmultiregimpl2_regs0 <= hdmi2usbsoc_hdmi_in0_edid_sda_i_async;
	xilinxmultiregimpl2_regs1 <= xilinxmultiregimpl2_regs0;
	xilinxmultiregimpl3_regs0 <= hdmi2usbsoc_hdmi_in0_locked_async;
	xilinxmultiregimpl3_regs1 <= xilinxmultiregimpl3_regs0;
	xilinxmultiregimpl4_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_done_toggle_i;
	xilinxmultiregimpl4_regs1 <= xilinxmultiregimpl4_regs0;
	xilinxmultiregimpl5_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_done_toggle_i;
	xilinxmultiregimpl5_regs1 <= xilinxmultiregimpl5_regs0;
	xilinxmultiregimpl12_regs0 <= {hdmi2usbsoc_hdmi_in0_s6datacapture0_too_early, hdmi2usbsoc_hdmi_in0_s6datacapture0_too_late};
	xilinxmultiregimpl12_regs1 <= xilinxmultiregimpl12_regs0;
	xilinxmultiregimpl14_regs0 <= hdmi2usbsoc_hdmi_in0_charsync0_synced;
	xilinxmultiregimpl14_regs1 <= xilinxmultiregimpl14_regs0;
	xilinxmultiregimpl15_regs0 <= hdmi2usbsoc_hdmi_in0_charsync0_word_sel;
	xilinxmultiregimpl15_regs1 <= xilinxmultiregimpl15_regs0;
	xilinxmultiregimpl16_regs0 <= hdmi2usbsoc_hdmi_in0_wer0_toggle_i;
	xilinxmultiregimpl16_regs1 <= xilinxmultiregimpl16_regs0;
	xilinxmultiregimpl17_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_done_toggle_i;
	xilinxmultiregimpl17_regs1 <= xilinxmultiregimpl17_regs0;
	xilinxmultiregimpl18_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_done_toggle_i;
	xilinxmultiregimpl18_regs1 <= xilinxmultiregimpl18_regs0;
	xilinxmultiregimpl25_regs0 <= {hdmi2usbsoc_hdmi_in0_s6datacapture1_too_early, hdmi2usbsoc_hdmi_in0_s6datacapture1_too_late};
	xilinxmultiregimpl25_regs1 <= xilinxmultiregimpl25_regs0;
	xilinxmultiregimpl27_regs0 <= hdmi2usbsoc_hdmi_in0_charsync1_synced;
	xilinxmultiregimpl27_regs1 <= xilinxmultiregimpl27_regs0;
	xilinxmultiregimpl28_regs0 <= hdmi2usbsoc_hdmi_in0_charsync1_word_sel;
	xilinxmultiregimpl28_regs1 <= xilinxmultiregimpl28_regs0;
	xilinxmultiregimpl29_regs0 <= hdmi2usbsoc_hdmi_in0_wer1_toggle_i;
	xilinxmultiregimpl29_regs1 <= xilinxmultiregimpl29_regs0;
	xilinxmultiregimpl30_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_done_toggle_i;
	xilinxmultiregimpl30_regs1 <= xilinxmultiregimpl30_regs0;
	xilinxmultiregimpl31_regs0 <= hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_done_toggle_i;
	xilinxmultiregimpl31_regs1 <= xilinxmultiregimpl31_regs0;
	xilinxmultiregimpl38_regs0 <= {hdmi2usbsoc_hdmi_in0_s6datacapture2_too_early, hdmi2usbsoc_hdmi_in0_s6datacapture2_too_late};
	xilinxmultiregimpl38_regs1 <= xilinxmultiregimpl38_regs0;
	xilinxmultiregimpl40_regs0 <= hdmi2usbsoc_hdmi_in0_charsync2_synced;
	xilinxmultiregimpl40_regs1 <= xilinxmultiregimpl40_regs0;
	xilinxmultiregimpl41_regs0 <= hdmi2usbsoc_hdmi_in0_charsync2_word_sel;
	xilinxmultiregimpl41_regs1 <= xilinxmultiregimpl41_regs0;
	xilinxmultiregimpl42_regs0 <= hdmi2usbsoc_hdmi_in0_wer2_toggle_i;
	xilinxmultiregimpl42_regs1 <= xilinxmultiregimpl42_regs0;
	xilinxmultiregimpl43_regs0 <= hdmi2usbsoc_hdmi_in0_chansync_chan_synced;
	xilinxmultiregimpl43_regs1 <= xilinxmultiregimpl43_regs0;
	xilinxmultiregimpl44_regs0 <= hdmi2usbsoc_hdmi_in0_resdetection_hcounter_st;
	xilinxmultiregimpl44_regs1 <= xilinxmultiregimpl44_regs0;
	xilinxmultiregimpl45_regs0 <= hdmi2usbsoc_hdmi_in0_resdetection_vcounter_st;
	xilinxmultiregimpl45_regs1 <= xilinxmultiregimpl45_regs0;
	xilinxmultiregimpl46_regs0 <= hdmi2usbsoc_hdmi_in0_frame_fifo_graycounter0_q;
	xilinxmultiregimpl46_regs1 <= xilinxmultiregimpl46_regs0;
	xilinxmultiregimpl48_regs0 <= hdmi2usbsoc_hdmi_in0_frame_pix_overflow;
	xilinxmultiregimpl48_regs1 <= xilinxmultiregimpl48_regs0;
	xilinxmultiregimpl50_regs0 <= hdmi2usbsoc_hdmi_in0_frame_overflow_reset_ack_toggle_i;
	xilinxmultiregimpl50_regs1 <= xilinxmultiregimpl50_regs0;
	xilinxmultiregimpl51_regs0 <= hdmi_in1_scl;
	xilinxmultiregimpl51_regs1 <= xilinxmultiregimpl51_regs0;
	xilinxmultiregimpl52_regs0 <= hdmi2usbsoc_hdmi_in1_edid_sda_i_async;
	xilinxmultiregimpl52_regs1 <= xilinxmultiregimpl52_regs0;
	xilinxmultiregimpl53_regs0 <= hdmi2usbsoc_hdmi_in1_locked_async;
	xilinxmultiregimpl53_regs1 <= xilinxmultiregimpl53_regs0;
	xilinxmultiregimpl54_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_done_toggle_i;
	xilinxmultiregimpl54_regs1 <= xilinxmultiregimpl54_regs0;
	xilinxmultiregimpl55_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_done_toggle_i;
	xilinxmultiregimpl55_regs1 <= xilinxmultiregimpl55_regs0;
	xilinxmultiregimpl62_regs0 <= {hdmi2usbsoc_hdmi_in1_s6datacapture0_too_early, hdmi2usbsoc_hdmi_in1_s6datacapture0_too_late};
	xilinxmultiregimpl62_regs1 <= xilinxmultiregimpl62_regs0;
	xilinxmultiregimpl64_regs0 <= hdmi2usbsoc_hdmi_in1_charsync0_synced;
	xilinxmultiregimpl64_regs1 <= xilinxmultiregimpl64_regs0;
	xilinxmultiregimpl65_regs0 <= hdmi2usbsoc_hdmi_in1_charsync0_word_sel;
	xilinxmultiregimpl65_regs1 <= xilinxmultiregimpl65_regs0;
	xilinxmultiregimpl66_regs0 <= hdmi2usbsoc_hdmi_in1_wer0_toggle_i;
	xilinxmultiregimpl66_regs1 <= xilinxmultiregimpl66_regs0;
	xilinxmultiregimpl67_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_done_toggle_i;
	xilinxmultiregimpl67_regs1 <= xilinxmultiregimpl67_regs0;
	xilinxmultiregimpl68_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_done_toggle_i;
	xilinxmultiregimpl68_regs1 <= xilinxmultiregimpl68_regs0;
	xilinxmultiregimpl75_regs0 <= {hdmi2usbsoc_hdmi_in1_s6datacapture1_too_early, hdmi2usbsoc_hdmi_in1_s6datacapture1_too_late};
	xilinxmultiregimpl75_regs1 <= xilinxmultiregimpl75_regs0;
	xilinxmultiregimpl77_regs0 <= hdmi2usbsoc_hdmi_in1_charsync1_synced;
	xilinxmultiregimpl77_regs1 <= xilinxmultiregimpl77_regs0;
	xilinxmultiregimpl78_regs0 <= hdmi2usbsoc_hdmi_in1_charsync1_word_sel;
	xilinxmultiregimpl78_regs1 <= xilinxmultiregimpl78_regs0;
	xilinxmultiregimpl79_regs0 <= hdmi2usbsoc_hdmi_in1_wer1_toggle_i;
	xilinxmultiregimpl79_regs1 <= xilinxmultiregimpl79_regs0;
	xilinxmultiregimpl80_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_done_toggle_i;
	xilinxmultiregimpl80_regs1 <= xilinxmultiregimpl80_regs0;
	xilinxmultiregimpl81_regs0 <= hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_done_toggle_i;
	xilinxmultiregimpl81_regs1 <= xilinxmultiregimpl81_regs0;
	xilinxmultiregimpl88_regs0 <= {hdmi2usbsoc_hdmi_in1_s6datacapture2_too_early, hdmi2usbsoc_hdmi_in1_s6datacapture2_too_late};
	xilinxmultiregimpl88_regs1 <= xilinxmultiregimpl88_regs0;
	xilinxmultiregimpl90_regs0 <= hdmi2usbsoc_hdmi_in1_charsync2_synced;
	xilinxmultiregimpl90_regs1 <= xilinxmultiregimpl90_regs0;
	xilinxmultiregimpl91_regs0 <= hdmi2usbsoc_hdmi_in1_charsync2_word_sel;
	xilinxmultiregimpl91_regs1 <= xilinxmultiregimpl91_regs0;
	xilinxmultiregimpl92_regs0 <= hdmi2usbsoc_hdmi_in1_wer2_toggle_i;
	xilinxmultiregimpl92_regs1 <= xilinxmultiregimpl92_regs0;
	xilinxmultiregimpl93_regs0 <= hdmi2usbsoc_hdmi_in1_chansync_chan_synced;
	xilinxmultiregimpl93_regs1 <= xilinxmultiregimpl93_regs0;
	xilinxmultiregimpl94_regs0 <= hdmi2usbsoc_hdmi_in1_resdetection_hcounter_st;
	xilinxmultiregimpl94_regs1 <= xilinxmultiregimpl94_regs0;
	xilinxmultiregimpl95_regs0 <= hdmi2usbsoc_hdmi_in1_resdetection_vcounter_st;
	xilinxmultiregimpl95_regs1 <= xilinxmultiregimpl95_regs0;
	xilinxmultiregimpl96_regs0 <= hdmi2usbsoc_hdmi_in1_frame_fifo_graycounter0_q;
	xilinxmultiregimpl96_regs1 <= xilinxmultiregimpl96_regs0;
	xilinxmultiregimpl98_regs0 <= hdmi2usbsoc_hdmi_in1_frame_pix_overflow;
	xilinxmultiregimpl98_regs1 <= xilinxmultiregimpl98_regs0;
	xilinxmultiregimpl100_regs0 <= hdmi2usbsoc_hdmi_in1_frame_overflow_reset_ack_toggle_i;
	xilinxmultiregimpl100_regs1 <= xilinxmultiregimpl100_regs0;
	xilinxmultiregimpl101_regs0 <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_graycounter0_q;
	xilinxmultiregimpl101_regs1 <= xilinxmultiregimpl101_regs0;
	xilinxmultiregimpl104_regs0 <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_graycounter1_q;
	xilinxmultiregimpl104_regs1 <= xilinxmultiregimpl104_regs0;
	xilinxmultiregimpl106_regs0 <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_graycounter1_q;
	xilinxmultiregimpl106_regs1 <= xilinxmultiregimpl106_regs0;
	xilinxmultiregimpl107_regs0 <= hdmi2usbsoc_hdmi_out0_core_underflow_enable_storage;
	xilinxmultiregimpl107_regs1 <= xilinxmultiregimpl107_regs0;
	xilinxmultiregimpl109_regs0 <= hdmi2usbsoc_hdmi_out0_driver_clocking_locked_async;
	xilinxmultiregimpl109_regs1 <= xilinxmultiregimpl109_regs0;
	xilinxmultiregimpl110_regs0 <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_graycounter2_q;
	xilinxmultiregimpl110_regs1 <= xilinxmultiregimpl110_regs0;
	xilinxmultiregimpl113_regs0 <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_graycounter3_q;
	xilinxmultiregimpl113_regs1 <= xilinxmultiregimpl113_regs0;
	xilinxmultiregimpl115_regs0 <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_graycounter1_q;
	xilinxmultiregimpl115_regs1 <= xilinxmultiregimpl115_regs0;
	xilinxmultiregimpl116_regs0 <= hdmi2usbsoc_hdmi_out1_core_underflow_enable_storage;
	xilinxmultiregimpl116_regs1 <= xilinxmultiregimpl116_regs0;
	xilinxmultiregimpl119_regs0 <= encoder_cdc_graycounter1_q;
	xilinxmultiregimpl119_regs1 <= xilinxmultiregimpl119_regs0;
end

always @(posedge usb_clk) begin
	encoder_streamer_fifo_graycounter1_q_binary <= encoder_streamer_fifo_graycounter1_q_next_binary;
	encoder_streamer_fifo_graycounter1_q <= encoder_streamer_fifo_graycounter1_q_next;
	if (usb_rst) begin
		encoder_streamer_fifo_graycounter1_q <= 3'd0;
		encoder_streamer_fifo_graycounter1_q_binary <= 3'd0;
	end
	xilinxmultiregimpl120_regs0 <= encoder_streamer_fifo_graycounter0_q;
	xilinxmultiregimpl120_regs1 <= xilinxmultiregimpl120_regs0;
end

lm32_cpu #(
	.eba_reset(32'h00000000)
) lm32_cpu (
	.D_ACK_I(hdmi2usbsoc_hdmi2usbsoc_dbus_ack),
	.D_DAT_I(hdmi2usbsoc_hdmi2usbsoc_dbus_dat_r),
	.D_ERR_I(hdmi2usbsoc_hdmi2usbsoc_dbus_err),
	.D_RTY_I(1'd0),
	.I_ACK_I(hdmi2usbsoc_hdmi2usbsoc_ibus_ack),
	.I_DAT_I(hdmi2usbsoc_hdmi2usbsoc_ibus_dat_r),
	.I_ERR_I(hdmi2usbsoc_hdmi2usbsoc_ibus_err),
	.I_RTY_I(1'd0),
	.clk_i(sys_clk),
	.interrupt(hdmi2usbsoc_hdmi2usbsoc_interrupt),
	.rst_i(sys_rst),
	.D_ADR_O(hdmi2usbsoc_hdmi2usbsoc_d_adr_o),
	.D_BTE_O(hdmi2usbsoc_hdmi2usbsoc_dbus_bte),
	.D_CTI_O(hdmi2usbsoc_hdmi2usbsoc_dbus_cti),
	.D_CYC_O(hdmi2usbsoc_hdmi2usbsoc_dbus_cyc),
	.D_DAT_O(hdmi2usbsoc_hdmi2usbsoc_dbus_dat_w),
	.D_SEL_O(hdmi2usbsoc_hdmi2usbsoc_dbus_sel),
	.D_STB_O(hdmi2usbsoc_hdmi2usbsoc_dbus_stb),
	.D_WE_O(hdmi2usbsoc_hdmi2usbsoc_dbus_we),
	.I_ADR_O(hdmi2usbsoc_hdmi2usbsoc_i_adr_o),
	.I_BTE_O(hdmi2usbsoc_hdmi2usbsoc_ibus_bte),
	.I_CTI_O(hdmi2usbsoc_hdmi2usbsoc_ibus_cti),
	.I_CYC_O(hdmi2usbsoc_hdmi2usbsoc_ibus_cyc),
	.I_DAT_O(hdmi2usbsoc_hdmi2usbsoc_ibus_dat_w),
	.I_SEL_O(hdmi2usbsoc_hdmi2usbsoc_ibus_sel),
	.I_STB_O(hdmi2usbsoc_hdmi2usbsoc_ibus_stb),
	.I_WE_O(hdmi2usbsoc_hdmi2usbsoc_ibus_we)
);

reg [31:0] mem[0:8191];
reg [12:0] memadr;
always @(posedge sys_clk) begin
	memadr <= hdmi2usbsoc_hdmi2usbsoc_rom_adr;
end

assign hdmi2usbsoc_hdmi2usbsoc_rom_dat_r = mem[memadr];

initial begin
	$readmemh("mem.init", mem);
end

reg [31:0] mem_1[0:4095];
reg [11:0] memadr_1;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_hdmi2usbsoc_sram_we[0])
		mem_1[hdmi2usbsoc_hdmi2usbsoc_sram_adr][7:0] <= hdmi2usbsoc_hdmi2usbsoc_sram_dat_w[7:0];
	if (hdmi2usbsoc_hdmi2usbsoc_sram_we[1])
		mem_1[hdmi2usbsoc_hdmi2usbsoc_sram_adr][15:8] <= hdmi2usbsoc_hdmi2usbsoc_sram_dat_w[15:8];
	if (hdmi2usbsoc_hdmi2usbsoc_sram_we[2])
		mem_1[hdmi2usbsoc_hdmi2usbsoc_sram_adr][23:16] <= hdmi2usbsoc_hdmi2usbsoc_sram_dat_w[23:16];
	if (hdmi2usbsoc_hdmi2usbsoc_sram_we[3])
		mem_1[hdmi2usbsoc_hdmi2usbsoc_sram_adr][31:24] <= hdmi2usbsoc_hdmi2usbsoc_sram_dat_w[31:24];
	memadr_1 <= hdmi2usbsoc_hdmi2usbsoc_sram_adr;
end

assign hdmi2usbsoc_hdmi2usbsoc_sram_dat_r = mem_1[memadr_1];

reg [9:0] storage[0:15];
reg [9:0] memdat;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_we)
		storage[hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_adr] <= hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_dat_w;
	memdat <= storage[hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_wrport_dat_r = memdat;
assign hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_rdport_dat_r = storage[hdmi2usbsoc_hdmi2usbsoc_uart_tx_fifo_rdport_adr];

reg [9:0] storage_1[0:15];
reg [9:0] memdat_1;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_we)
		storage_1[hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_adr] <= hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_dat_w;
	memdat_1 <= storage_1[hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_wrport_dat_r = memdat_1;
assign hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_rdport_dat_r = storage_1[hdmi2usbsoc_hdmi2usbsoc_uart_rx_fifo_rdport_adr];

reg [7:0] mem_2[0:11];
reg [3:0] memadr_2;
always @(posedge sys_clk) begin
	memadr_2 <= hdmi2usbsoc_sram2_adr;
end

assign hdmi2usbsoc_sram2_dat_r = mem_2[memadr_2];

initial begin
	$readmemh("mem_2.init", mem_2);
end

IBUFG IBUFG(
	.I(clk100),
	.O(hdmi2usbsoc_crg_clk100a)
);

BUFIO2 #(
	.DIVIDE(1'd1),
	.DIVIDE_BYPASS("TRUE"),
	.I_INVERT("FALSE")
) BUFIO2 (
	.I(hdmi2usbsoc_crg_clk100a),
	.DIVCLK(hdmi2usbsoc_crg_clk100b)
);

PLL_ADV #(
	.BANDWIDTH("OPTIMIZED"),
	.CLKFBOUT_MULT(3'd6),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(10.0),
	.CLKIN2_PERIOD(0.0),
	.CLKOUT0_DIVIDE(2'd2),
	.CLKOUT0_DUTY_CYCLE(0.5),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(4'd9),
	.CLKOUT1_DUTY_CYCLE(0.5),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(3'd4),
	.CLKOUT2_DUTY_CYCLE(0.5),
	.CLKOUT2_PHASE(270.0),
	.CLKOUT3_DIVIDE(3'd4),
	.CLKOUT3_DUTY_CYCLE(0.5),
	.CLKOUT3_PHASE(250.0),
	.CLKOUT4_DIVIDE(4'd12),
	.CLKOUT4_DUTY_CYCLE(0.5),
	.CLKOUT4_PHASE(0.0),
	.CLKOUT5_DIVIDE(4'd8),
	.CLKOUT5_DUTY_CYCLE(0.5),
	.CLKOUT5_PHASE(0.0),
	.CLK_FEEDBACK("CLKFBOUT"),
	.COMPENSATION("INTERNAL"),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER(0.01),
	.SIM_DEVICE("SPARTAN6")
) crg_pll_adv (
	.CLKFBIN(hdmi2usbsoc_crg_pll_fb),
	.CLKIN1(hdmi2usbsoc_crg_clk100b),
	.CLKIN2(1'd0),
	.CLKINSEL(1'd1),
	.DADDR(1'd0),
	.DCLK(1'd0),
	.DEN(1'd0),
	.DI(1'd0),
	.DWE(1'd0),
	.REL(1'd0),
	.RST(1'd0),
	.CLKFBOUT(hdmi2usbsoc_crg_pll_fb),
	.CLKOUT0(hdmi2usbsoc_crg_unbuf_sdram_full),
	.CLKOUT1(hdmi2usbsoc_crg_unbuf_encoder),
	.CLKOUT2(hdmi2usbsoc_crg_unbuf_sdram_half_a),
	.CLKOUT3(hdmi2usbsoc_crg_unbuf_sdram_half_b),
	.CLKOUT4(hdmi2usbsoc_crg_unbuf_unused),
	.CLKOUT5(hdmi2usbsoc_crg_unbuf_sys),
	.LOCKED(hdmi2usbsoc_crg_pll_lckd)
);

BUFG sys_bufg(
	.I(hdmi2usbsoc_crg_unbuf_sys),
	.O(sys_clk)
);

BUFPLL #(
	.DIVIDE(3'd4)
) sdram_full_bufpll (
	.GCLK(sys_clk),
	.LOCKED(hdmi2usbsoc_crg_pll_lckd),
	.PLLIN(hdmi2usbsoc_crg_unbuf_sdram_full),
	.IOCLK(sdram_full_wr_clk),
	.SERDESSTROBE(hdmi2usbsoc_crg_clk4x_wr_strb)
);

BUFG sdram_half_a_bufpll(
	.I(hdmi2usbsoc_crg_unbuf_sdram_half_a),
	.O(sdram_half_clk)
);

BUFG sdram_half_b_bufpll(
	.I(hdmi2usbsoc_crg_unbuf_sdram_half_b),
	.O(hdmi2usbsoc_crg_clk_sdram_half_shifted)
);

ODDR2 #(
	.DDR_ALIGNMENT("NONE"),
	.INIT(1'd0),
	.SRTYPE("SYNC")
) ODDR2 (
	.C0(hdmi2usbsoc_crg_clk_sdram_half_shifted),
	.C1((~hdmi2usbsoc_crg_clk_sdram_half_shifted)),
	.CE(1'd1),
	.D0(1'd1),
	.D1(1'd0),
	.R(1'd0),
	.S(1'd0),
	.Q(hdmi2usbsoc_crg_output_clk)
);

OBUFDS OBUFDS(
	.I(hdmi2usbsoc_crg_output_clk),
	.O(ddram_clock_p),
	.OB(ddram_clock_n)
);

DCM_CLKGEN #(
	.CLKFXDV_DIVIDE(2'd2),
	.CLKFX_DIVIDE(3'd4),
	.CLKFX_MD_MAX(0.5),
	.CLKFX_MULTIPLY(2'd2),
	.CLKIN_PERIOD(10.0),
	.SPREAD_SPECTRUM("NONE"),
	.STARTUP_WAIT("FALSE")
) crg_periph_dcm_clkgen (
	.CLKIN(hdmi2usbsoc_crg_clk100a),
	.FREEZEDCM(1'd0),
	.RST(sys_rst),
	.CLKFX(base50_clk),
	.LOCKED(hdmi2usbsoc_crg_dcm_base50_locked)
);

BUFG encoder_bufg(
	.I(hdmi2usbsoc_crg_unbuf_encoder),
	.O(encoder_clk)
);

DNA_PORT DNA_PORT(
	.CLK(hdmi2usbsoc_dna_cnt[0]),
	.DIN(hdmi2usbsoc_dna_status[56]),
	.READ((hdmi2usbsoc_dna_cnt < 2'd2)),
	.SHIFT(1'd1),
	.DOUT(hdmi2usbsoc_dna_do)
);

assign spiflash4x_dq = hdmi2usbsoc_oe ? hdmi2usbsoc_o : 4'bz;
assign hdmi2usbsoc_i0 = spiflash4x_dq;

ODDR2 #(
	.DDR_ALIGNMENT("C0"),
	.INIT(1'd0),
	.SRTYPE("ASYNC")
) ODDR2_1 (
	.C0(sdram_half_clk),
	.C1(hdmi2usbsoc_ddrphy_sdram_half_clk_n),
	.CE(1'd1),
	.D0(1'd0),
	.D1(1'd1),
	.R(1'd0),
	.S(1'd0),
	.Q(hdmi2usbsoc_ddrphy_dqs_o[0])
);

ODDR2 #(
	.DDR_ALIGNMENT("C0"),
	.INIT(1'd0),
	.SRTYPE("ASYNC")
) ODDR2_2 (
	.C0(sdram_half_clk),
	.C1(hdmi2usbsoc_ddrphy_sdram_half_clk_n),
	.CE(1'd1),
	.D0(hdmi2usbsoc_ddrphy_dqs_t_d0),
	.D1(hdmi2usbsoc_ddrphy_dqs_t_d1),
	.R(1'd0),
	.S(1'd0),
	.Q(hdmi2usbsoc_ddrphy_dqs_t[0])
);

OBUFTDS OBUFTDS(
	.I(hdmi2usbsoc_ddrphy_dqs_o[0]),
	.T(hdmi2usbsoc_ddrphy_dqs_t[0]),
	.O(ddram_dqs[0]),
	.OB(ddram_dqs_n[0])
);

ODDR2 #(
	.DDR_ALIGNMENT("C0"),
	.INIT(1'd0),
	.SRTYPE("ASYNC")
) ODDR2_3 (
	.C0(sdram_half_clk),
	.C1(hdmi2usbsoc_ddrphy_sdram_half_clk_n),
	.CE(1'd1),
	.D0(1'd0),
	.D1(1'd1),
	.R(1'd0),
	.S(1'd0),
	.Q(hdmi2usbsoc_ddrphy_dqs_o[1])
);

ODDR2 #(
	.DDR_ALIGNMENT("C0"),
	.INIT(1'd0),
	.SRTYPE("ASYNC")
) ODDR2_4 (
	.C0(sdram_half_clk),
	.C1(hdmi2usbsoc_ddrphy_sdram_half_clk_n),
	.CE(1'd1),
	.D0(hdmi2usbsoc_ddrphy_dqs_t_d0),
	.D1(hdmi2usbsoc_ddrphy_dqs_t_d1),
	.R(1'd0),
	.S(1'd0),
	.Q(hdmi2usbsoc_ddrphy_dqs_t[1])
);

OBUFTDS OBUFTDS_1(
	.I(hdmi2usbsoc_ddrphy_dqs_o[1]),
	.T(hdmi2usbsoc_ddrphy_dqs_t[1]),
	.O(ddram_dqs[1]),
	.OB(ddram_dqs_n[1])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy0[0]),
	.D2(slice_proxy1[0]),
	.D3(slice_proxy2[0]),
	.D4(slice_proxy3[0]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[0]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[0])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[0]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[16]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[0]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[16]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[0])
);

IOBUF IOBUF(
	.I(hdmi2usbsoc_ddrphy_dq_o[0]),
	.T(hdmi2usbsoc_ddrphy_dq_t[0]),
	.IO(ddram_dq[0]),
	.O(hdmi2usbsoc_ddrphy_dq_i[0])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_1 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy4[1]),
	.D2(slice_proxy5[1]),
	.D3(slice_proxy6[1]),
	.D4(slice_proxy7[1]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[1]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[1])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_1 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[1]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[17]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[1]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[17]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[1])
);

IOBUF IOBUF_1(
	.I(hdmi2usbsoc_ddrphy_dq_o[1]),
	.T(hdmi2usbsoc_ddrphy_dq_t[1]),
	.IO(ddram_dq[1]),
	.O(hdmi2usbsoc_ddrphy_dq_i[1])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_2 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy8[2]),
	.D2(slice_proxy9[2]),
	.D3(slice_proxy10[2]),
	.D4(slice_proxy11[2]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[2]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[2])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_2 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[2]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[18]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[2]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[18]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[2])
);

IOBUF IOBUF_2(
	.I(hdmi2usbsoc_ddrphy_dq_o[2]),
	.T(hdmi2usbsoc_ddrphy_dq_t[2]),
	.IO(ddram_dq[2]),
	.O(hdmi2usbsoc_ddrphy_dq_i[2])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_3 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy12[3]),
	.D2(slice_proxy13[3]),
	.D3(slice_proxy14[3]),
	.D4(slice_proxy15[3]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[3]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[3])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_3 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[3]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[19]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[3]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[19]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[3])
);

IOBUF IOBUF_3(
	.I(hdmi2usbsoc_ddrphy_dq_o[3]),
	.T(hdmi2usbsoc_ddrphy_dq_t[3]),
	.IO(ddram_dq[3]),
	.O(hdmi2usbsoc_ddrphy_dq_i[3])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_4 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy16[4]),
	.D2(slice_proxy17[4]),
	.D3(slice_proxy18[4]),
	.D4(slice_proxy19[4]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[4]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[4])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_4 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[4]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[20]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[4]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[20]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[4])
);

IOBUF IOBUF_4(
	.I(hdmi2usbsoc_ddrphy_dq_o[4]),
	.T(hdmi2usbsoc_ddrphy_dq_t[4]),
	.IO(ddram_dq[4]),
	.O(hdmi2usbsoc_ddrphy_dq_i[4])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_5 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy20[5]),
	.D2(slice_proxy21[5]),
	.D3(slice_proxy22[5]),
	.D4(slice_proxy23[5]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[5]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[5])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_5 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[5]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[21]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[5]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[21]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[5])
);

IOBUF IOBUF_5(
	.I(hdmi2usbsoc_ddrphy_dq_o[5]),
	.T(hdmi2usbsoc_ddrphy_dq_t[5]),
	.IO(ddram_dq[5]),
	.O(hdmi2usbsoc_ddrphy_dq_i[5])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_6 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy24[6]),
	.D2(slice_proxy25[6]),
	.D3(slice_proxy26[6]),
	.D4(slice_proxy27[6]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[6]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[6])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_6 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[6]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[22]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[6]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[22]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[6])
);

IOBUF IOBUF_6(
	.I(hdmi2usbsoc_ddrphy_dq_o[6]),
	.T(hdmi2usbsoc_ddrphy_dq_t[6]),
	.IO(ddram_dq[6]),
	.O(hdmi2usbsoc_ddrphy_dq_i[6])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_7 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy28[7]),
	.D2(slice_proxy29[7]),
	.D3(slice_proxy30[7]),
	.D4(slice_proxy31[7]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[7]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[7])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_7 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[7]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[23]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[7]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[23]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[7])
);

IOBUF IOBUF_7(
	.I(hdmi2usbsoc_ddrphy_dq_o[7]),
	.T(hdmi2usbsoc_ddrphy_dq_t[7]),
	.IO(ddram_dq[7]),
	.O(hdmi2usbsoc_ddrphy_dq_i[7])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_8 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy32[8]),
	.D2(slice_proxy33[8]),
	.D3(slice_proxy34[8]),
	.D4(slice_proxy35[8]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[8]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[8])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_8 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[8]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[24]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[8]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[24]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[8])
);

IOBUF IOBUF_8(
	.I(hdmi2usbsoc_ddrphy_dq_o[8]),
	.T(hdmi2usbsoc_ddrphy_dq_t[8]),
	.IO(ddram_dq[8]),
	.O(hdmi2usbsoc_ddrphy_dq_i[8])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_9 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy36[9]),
	.D2(slice_proxy37[9]),
	.D3(slice_proxy38[9]),
	.D4(slice_proxy39[9]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[9]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[9])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_9 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[9]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[25]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[9]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[25]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[9])
);

IOBUF IOBUF_9(
	.I(hdmi2usbsoc_ddrphy_dq_o[9]),
	.T(hdmi2usbsoc_ddrphy_dq_t[9]),
	.IO(ddram_dq[9]),
	.O(hdmi2usbsoc_ddrphy_dq_i[9])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_10 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy40[10]),
	.D2(slice_proxy41[10]),
	.D3(slice_proxy42[10]),
	.D4(slice_proxy43[10]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[10]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[10])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_10 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[10]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[26]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[10]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[26]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[10])
);

IOBUF IOBUF_10(
	.I(hdmi2usbsoc_ddrphy_dq_o[10]),
	.T(hdmi2usbsoc_ddrphy_dq_t[10]),
	.IO(ddram_dq[10]),
	.O(hdmi2usbsoc_ddrphy_dq_i[10])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_11 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy44[11]),
	.D2(slice_proxy45[11]),
	.D3(slice_proxy46[11]),
	.D4(slice_proxy47[11]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[11]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[11])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_11 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[11]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[27]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[11]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[27]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[11])
);

IOBUF IOBUF_11(
	.I(hdmi2usbsoc_ddrphy_dq_o[11]),
	.T(hdmi2usbsoc_ddrphy_dq_t[11]),
	.IO(ddram_dq[11]),
	.O(hdmi2usbsoc_ddrphy_dq_i[11])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_12 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy48[12]),
	.D2(slice_proxy49[12]),
	.D3(slice_proxy50[12]),
	.D4(slice_proxy51[12]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[12]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[12])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_12 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[12]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[28]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[12]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[28]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[12])
);

IOBUF IOBUF_12(
	.I(hdmi2usbsoc_ddrphy_dq_o[12]),
	.T(hdmi2usbsoc_ddrphy_dq_t[12]),
	.IO(ddram_dq[12]),
	.O(hdmi2usbsoc_ddrphy_dq_i[12])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_13 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy52[13]),
	.D2(slice_proxy53[13]),
	.D3(slice_proxy54[13]),
	.D4(slice_proxy55[13]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[13]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[13])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_13 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[13]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[29]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[13]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[29]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[13])
);

IOBUF IOBUF_13(
	.I(hdmi2usbsoc_ddrphy_dq_o[13]),
	.T(hdmi2usbsoc_ddrphy_dq_t[13]),
	.IO(ddram_dq[13]),
	.O(hdmi2usbsoc_ddrphy_dq_i[13])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_14 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy56[14]),
	.D2(slice_proxy57[14]),
	.D3(slice_proxy58[14]),
	.D4(slice_proxy59[14]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[14]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[14])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_14 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[14]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[30]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[14]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[30]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[14])
);

IOBUF IOBUF_14(
	.I(hdmi2usbsoc_ddrphy_dq_o[14]),
	.T(hdmi2usbsoc_ddrphy_dq_t[14]),
	.IO(ddram_dq[14]),
	.O(hdmi2usbsoc_ddrphy_dq_i[14])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_15 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy60[15]),
	.D2(slice_proxy61[15]),
	.D3(slice_proxy62[15]),
	.D4(slice_proxy63[15]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.T1(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T2(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T3(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.T4(hdmi2usbsoc_ddrphy_drive_dq_n1),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_ddrphy_dq_o[15]),
	.TQ(hdmi2usbsoc_ddrphy_dq_t[15])
);

ISERDES2 #(
	.BITSLIP_ENABLE("TRUE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd4),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("NONE")
) ISERDES2_15 (
	.BITSLIP(hdmi2usbsoc_ddrphy_bitslip_inc),
	.CE0(1'd1),
	.CLK0(sdram_full_rd_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D(hdmi2usbsoc_ddrphy_dq_i[15]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_rd_strb),
	.RST(sys_rst),
	.Q1(hdmi2usbsoc_ddrphy_record0_rddata[31]),
	.Q2(hdmi2usbsoc_ddrphy_record0_rddata[15]),
	.Q3(hdmi2usbsoc_ddrphy_record1_rddata[31]),
	.Q4(hdmi2usbsoc_ddrphy_record1_rddata[15])
);

IOBUF IOBUF_15(
	.I(hdmi2usbsoc_ddrphy_dq_o[15]),
	.T(hdmi2usbsoc_ddrphy_dq_t[15]),
	.IO(ddram_dq[15]),
	.O(hdmi2usbsoc_ddrphy_dq_i[15])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_16 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy64[0]),
	.D2(slice_proxy65[0]),
	.D3(slice_proxy66[0]),
	.D4(slice_proxy67[0]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.TCE(1'd0),
	.TRAIN(1'd0),
	.OQ(ddram_dm[0])
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd4),
	.OUTPUT_MODE("SINGLE_ENDED"),
	.SERDES_MODE("NONE")
) OSERDES2_17 (
	.CLK0(sdram_full_wr_clk),
	.CLK1(1'd0),
	.CLKDIV(sys_clk),
	.D1(slice_proxy68[1]),
	.D2(slice_proxy69[1]),
	.D3(slice_proxy70[1]),
	.D4(slice_proxy71[1]),
	.IOCE(hdmi2usbsoc_ddrphy_clk4x_wr_strb),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.SHIFTIN3(1'd0),
	.SHIFTIN4(1'd0),
	.TCE(1'd0),
	.TRAIN(1'd0),
	.OQ(ddram_dm[1])
);

reg [23:0] storage_2[0:7];
reg [23:0] memdat_2;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine0_wrport_we)
		storage_2[hdmi2usbsoc_sdram_bankmachine0_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine0_wrport_dat_w;
	memdat_2 <= storage_2[hdmi2usbsoc_sdram_bankmachine0_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine0_wrport_dat_r = memdat_2;
assign hdmi2usbsoc_sdram_bankmachine0_rdport_dat_r = storage_2[hdmi2usbsoc_sdram_bankmachine0_rdport_adr];

reg [23:0] storage_3[0:7];
reg [23:0] memdat_3;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine1_wrport_we)
		storage_3[hdmi2usbsoc_sdram_bankmachine1_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine1_wrport_dat_w;
	memdat_3 <= storage_3[hdmi2usbsoc_sdram_bankmachine1_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine1_wrport_dat_r = memdat_3;
assign hdmi2usbsoc_sdram_bankmachine1_rdport_dat_r = storage_3[hdmi2usbsoc_sdram_bankmachine1_rdport_adr];

reg [23:0] storage_4[0:7];
reg [23:0] memdat_4;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine2_wrport_we)
		storage_4[hdmi2usbsoc_sdram_bankmachine2_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine2_wrport_dat_w;
	memdat_4 <= storage_4[hdmi2usbsoc_sdram_bankmachine2_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine2_wrport_dat_r = memdat_4;
assign hdmi2usbsoc_sdram_bankmachine2_rdport_dat_r = storage_4[hdmi2usbsoc_sdram_bankmachine2_rdport_adr];

reg [23:0] storage_5[0:7];
reg [23:0] memdat_5;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine3_wrport_we)
		storage_5[hdmi2usbsoc_sdram_bankmachine3_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine3_wrport_dat_w;
	memdat_5 <= storage_5[hdmi2usbsoc_sdram_bankmachine3_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine3_wrport_dat_r = memdat_5;
assign hdmi2usbsoc_sdram_bankmachine3_rdport_dat_r = storage_5[hdmi2usbsoc_sdram_bankmachine3_rdport_adr];

reg [23:0] storage_6[0:7];
reg [23:0] memdat_6;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine4_wrport_we)
		storage_6[hdmi2usbsoc_sdram_bankmachine4_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine4_wrport_dat_w;
	memdat_6 <= storage_6[hdmi2usbsoc_sdram_bankmachine4_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine4_wrport_dat_r = memdat_6;
assign hdmi2usbsoc_sdram_bankmachine4_rdport_dat_r = storage_6[hdmi2usbsoc_sdram_bankmachine4_rdport_adr];

reg [23:0] storage_7[0:7];
reg [23:0] memdat_7;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine5_wrport_we)
		storage_7[hdmi2usbsoc_sdram_bankmachine5_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine5_wrport_dat_w;
	memdat_7 <= storage_7[hdmi2usbsoc_sdram_bankmachine5_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine5_wrport_dat_r = memdat_7;
assign hdmi2usbsoc_sdram_bankmachine5_rdport_dat_r = storage_7[hdmi2usbsoc_sdram_bankmachine5_rdport_adr];

reg [23:0] storage_8[0:7];
reg [23:0] memdat_8;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine6_wrport_we)
		storage_8[hdmi2usbsoc_sdram_bankmachine6_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine6_wrport_dat_w;
	memdat_8 <= storage_8[hdmi2usbsoc_sdram_bankmachine6_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine6_wrport_dat_r = memdat_8;
assign hdmi2usbsoc_sdram_bankmachine6_rdport_dat_r = storage_8[hdmi2usbsoc_sdram_bankmachine6_rdport_adr];

reg [23:0] storage_9[0:7];
reg [23:0] memdat_9;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sdram_bankmachine7_wrport_we)
		storage_9[hdmi2usbsoc_sdram_bankmachine7_wrport_adr] <= hdmi2usbsoc_sdram_bankmachine7_wrport_dat_w;
	memdat_9 <= storage_9[hdmi2usbsoc_sdram_bankmachine7_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_sdram_bankmachine7_wrport_dat_r = memdat_9;
assign hdmi2usbsoc_sdram_bankmachine7_rdport_dat_r = storage_9[hdmi2usbsoc_sdram_bankmachine7_rdport_adr];

reg [63:0] data_mem[0:1023];
reg [9:0] memadr_3;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_data_port_we[0])
		data_mem[hdmi2usbsoc_data_port_adr][7:0] <= hdmi2usbsoc_data_port_dat_w[7:0];
	if (hdmi2usbsoc_data_port_we[1])
		data_mem[hdmi2usbsoc_data_port_adr][15:8] <= hdmi2usbsoc_data_port_dat_w[15:8];
	if (hdmi2usbsoc_data_port_we[2])
		data_mem[hdmi2usbsoc_data_port_adr][23:16] <= hdmi2usbsoc_data_port_dat_w[23:16];
	if (hdmi2usbsoc_data_port_we[3])
		data_mem[hdmi2usbsoc_data_port_adr][31:24] <= hdmi2usbsoc_data_port_dat_w[31:24];
	if (hdmi2usbsoc_data_port_we[4])
		data_mem[hdmi2usbsoc_data_port_adr][39:32] <= hdmi2usbsoc_data_port_dat_w[39:32];
	if (hdmi2usbsoc_data_port_we[5])
		data_mem[hdmi2usbsoc_data_port_adr][47:40] <= hdmi2usbsoc_data_port_dat_w[47:40];
	if (hdmi2usbsoc_data_port_we[6])
		data_mem[hdmi2usbsoc_data_port_adr][55:48] <= hdmi2usbsoc_data_port_dat_w[55:48];
	if (hdmi2usbsoc_data_port_we[7])
		data_mem[hdmi2usbsoc_data_port_adr][63:56] <= hdmi2usbsoc_data_port_dat_w[63:56];
	memadr_3 <= hdmi2usbsoc_data_port_adr;
end

assign hdmi2usbsoc_data_port_dat_r = data_mem[memadr_3];

reg [21:0] tag_mem[0:1023];
reg [9:0] memadr_4;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_tag_port_we)
		tag_mem[hdmi2usbsoc_tag_port_adr] <= hdmi2usbsoc_tag_port_dat_w;
	memadr_4 <= hdmi2usbsoc_tag_port_adr;
end

assign hdmi2usbsoc_tag_port_dat_r = tag_mem[memadr_4];

reg [7:0] edid_mem[0:127];
reg [6:0] memadr_5;
reg [6:0] memadr_6;
always @(posedge sys_clk) begin
	memadr_5 <= hdmi2usbsoc_hdmi_in0_edid_adr;
end

always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sram0_we)
		edid_mem[hdmi2usbsoc_sram0_adr] <= hdmi2usbsoc_sram0_dat_w;
	memadr_6 <= hdmi2usbsoc_sram0_adr;
end

assign hdmi2usbsoc_hdmi_in0_edid_dat_r = edid_mem[memadr_5];
assign hdmi2usbsoc_sram0_dat_r = edid_mem[memadr_6];

initial begin
	$readmemh("edid_mem.init", edid_mem);
end

assign hdmi_in0_sda = hdmi2usbsoc_hdmi_in0_edid_sda_drv_reg ? 1'd0 : 1'bz;
assign hdmi2usbsoc_hdmi_in0_edid_sda_i_async = hdmi_in0_sda;

IBUFDS hdmi_in_ibufds(
	.I(hdmi_in0_clk_p),
	.IB(hdmi_in0_clk_n),
	.O(hdmi2usbsoc_hdmi_in0_clk_input)
);

PLL_ADV #(
	.CLKFBOUT_MULT(4'd10),
	.CLKOUT0_DIVIDE(1'd1),
	.CLKOUT1_DIVIDE(3'd5),
	.CLKOUT2_DIVIDE(4'd10),
	.COMPENSATION("INTERNAL")
) hdmi_in_pll_adv (
	.CLKFBIN(hdmi2usbsoc_hdmi_in0_clkfbout),
	.CLKIN1(hdmi2usbsoc_hdmi_in0_clk_input),
	.CLKINSEL(1'd1),
	.DADDR(hdmi2usbsoc_hdmi_in0_pll_adr_storage),
	.DCLK(sys_clk),
	.DEN((hdmi2usbsoc_hdmi_in0_pll_read_re | hdmi2usbsoc_hdmi_in0_pll_write_re)),
	.DI(hdmi2usbsoc_hdmi_in0_pll_dat_w_storage),
	.DWE(hdmi2usbsoc_hdmi_in0_pll_write_re),
	.RST(hdmi2usbsoc_hdmi_in0_pll_reset_storage),
	.CLKFBOUT(hdmi2usbsoc_hdmi_in0_clkfbout),
	.CLKOUT0(hdmi2usbsoc_hdmi_in0_pll_clk0),
	.CLKOUT1(hdmi2usbsoc_hdmi_in0_pll_clk1),
	.CLKOUT2(hdmi2usbsoc_hdmi_in0_pll_clk2),
	.DO(hdmi2usbsoc_hdmi_in0_pll_dat_r_status),
	.DRDY(hdmi2usbsoc_hdmi_in0_pll_drdy),
	.LOCKED(hdmi2usbsoc_hdmi_in0_pll_locked)
);

BUFPLL #(
	.DIVIDE(3'd5)
) hdmi_in_bufpll (
	.GCLK(hdmi_in0_pix2x_clk),
	.LOCKED(hdmi2usbsoc_hdmi_in0_pll_locked),
	.PLLIN(hdmi2usbsoc_hdmi_in0_pll_clk0),
	.IOCLK(hdmi_in0_pix10x_clk),
	.LOCK(hdmi2usbsoc_hdmi_in0_locked_async),
	.SERDESSTROBE(hdmi2usbsoc_hdmi_in0_serdesstrobe)
);

BUFG hdmi_in_pix2x_bufg(
	.I(hdmi2usbsoc_hdmi_in0_pll_clk1),
	.O(hdmi_in0_pix2x_clk)
);

BUFG hdmi_in_pix_bufg(
	.I(hdmi2usbsoc_hdmi_in0_pll_clk2),
	.O(hdmi_in0_pix_clk)
);

IBUFDS IBUFDS(
	.I(hdmi_in0_data0_p),
	.IB(hdmi_in0_data0_n),
	.O(hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_se)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("STAY_AT_LIMIT"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("MASTER")
) IODELAY2 (
	.CAL(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_cal),
	.CE(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_ce),
	.CLK(hdmi_in0_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_se),
	.INC(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_inc),
	.IOCLK0(hdmi_in0_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_master_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_delayed_master)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("WRAPAROUND"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("SLAVE")
) IODELAY2_1 (
	.CAL(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_cal),
	.CE(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_ce),
	.CLK(hdmi_in0_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_se),
	.INC(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_inc),
	.IOCLK0(hdmi_in0_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in0_s6datacapture0_delay_slave_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_delayed_slave)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("MASTER")
) ISERDES2_16 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in0_pix10x_clk),
	.CLKDIV(hdmi_in0_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_delayed_master),
	.IOCE(hdmi2usbsoc_hdmi_in0_s6datacapture0_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_edge),
	.INCDEC(hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_incdec),
	.Q1(hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr2[1]),
	.Q2(hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr2[2]),
	.Q3(hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr2[3]),
	.Q4(hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr2[4]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_cascade),
	.VALID(hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_valid)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("SLAVE")
) ISERDES2_17 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in0_pix10x_clk),
	.CLKDIV(hdmi_in0_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in0_s6datacapture0_pad_delayed_slave),
	.IOCE(hdmi2usbsoc_hdmi_in0_s6datacapture0_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_cascade),
	.Q4(hdmi2usbsoc_hdmi_in0_s6datacapture0_dsr2[0]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in0_s6datacapture0_pd_edge)
);

IBUFDS IBUFDS_1(
	.I(hdmi_in0_data1_p),
	.IB(hdmi_in0_data1_n),
	.O(hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_se)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("STAY_AT_LIMIT"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("MASTER")
) IODELAY2_2 (
	.CAL(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_cal),
	.CE(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_ce),
	.CLK(hdmi_in0_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_se),
	.INC(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_inc),
	.IOCLK0(hdmi_in0_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_master_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_delayed_master)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("WRAPAROUND"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("SLAVE")
) IODELAY2_3 (
	.CAL(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_cal),
	.CE(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_ce),
	.CLK(hdmi_in0_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_se),
	.INC(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_inc),
	.IOCLK0(hdmi_in0_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in0_s6datacapture1_delay_slave_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_delayed_slave)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("MASTER")
) ISERDES2_18 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in0_pix10x_clk),
	.CLKDIV(hdmi_in0_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_delayed_master),
	.IOCE(hdmi2usbsoc_hdmi_in0_s6datacapture1_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_edge),
	.INCDEC(hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_incdec),
	.Q1(hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr2[1]),
	.Q2(hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr2[2]),
	.Q3(hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr2[3]),
	.Q4(hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr2[4]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_cascade),
	.VALID(hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_valid)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("SLAVE")
) ISERDES2_19 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in0_pix10x_clk),
	.CLKDIV(hdmi_in0_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in0_s6datacapture1_pad_delayed_slave),
	.IOCE(hdmi2usbsoc_hdmi_in0_s6datacapture1_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_cascade),
	.Q4(hdmi2usbsoc_hdmi_in0_s6datacapture1_dsr2[0]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in0_s6datacapture1_pd_edge)
);

IBUFDS IBUFDS_2(
	.I(hdmi_in0_data2_p),
	.IB(hdmi_in0_data2_n),
	.O(hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_se)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("STAY_AT_LIMIT"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("MASTER")
) IODELAY2_4 (
	.CAL(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_cal),
	.CE(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_ce),
	.CLK(hdmi_in0_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_se),
	.INC(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_inc),
	.IOCLK0(hdmi_in0_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_master_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_delayed_master)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("WRAPAROUND"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("SLAVE")
) IODELAY2_5 (
	.CAL(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_cal),
	.CE(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_ce),
	.CLK(hdmi_in0_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_se),
	.INC(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_inc),
	.IOCLK0(hdmi_in0_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in0_s6datacapture2_delay_slave_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_delayed_slave)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("MASTER")
) ISERDES2_20 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in0_pix10x_clk),
	.CLKDIV(hdmi_in0_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_delayed_master),
	.IOCE(hdmi2usbsoc_hdmi_in0_s6datacapture2_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_edge),
	.INCDEC(hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_incdec),
	.Q1(hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr2[1]),
	.Q2(hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr2[2]),
	.Q3(hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr2[3]),
	.Q4(hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr2[4]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_cascade),
	.VALID(hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_valid)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("SLAVE")
) ISERDES2_21 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in0_pix10x_clk),
	.CLKDIV(hdmi_in0_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in0_s6datacapture2_pad_delayed_slave),
	.IOCE(hdmi2usbsoc_hdmi_in0_s6datacapture2_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_cascade),
	.Q4(hdmi2usbsoc_hdmi_in0_s6datacapture2_dsr2[0]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in0_s6datacapture2_pd_edge)
);

reg [20:0] storage_10[0:7];
reg [2:0] memadr_7;
always @(posedge hdmi_in0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_we)
		storage_10[hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_adr] <= hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_w;
	memadr_7 <= hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_wrport_dat_r = storage_10[memadr_7];
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_rdport_dat_r = storage_10[hdmi2usbsoc_hdmi_in0_chansync_syncbuffer0_rdport_adr];

reg [20:0] storage_11[0:7];
reg [2:0] memadr_8;
always @(posedge hdmi_in0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_we)
		storage_11[hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_adr] <= hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_w;
	memadr_8 <= hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_wrport_dat_r = storage_11[memadr_8];
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_rdport_dat_r = storage_11[hdmi2usbsoc_hdmi_in0_chansync_syncbuffer1_rdport_adr];

reg [20:0] storage_12[0:7];
reg [2:0] memadr_9;
always @(posedge hdmi_in0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_we)
		storage_12[hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_adr] <= hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_w;
	memadr_9 <= hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_wrport_dat_r = storage_12[memadr_9];
assign hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_rdport_dat_r = storage_12[hdmi2usbsoc_hdmi_in0_chansync_syncbuffer2_rdport_adr];

reg [66:0] storage_13[0:511];
reg [8:0] memadr_10;
reg [8:0] memadr_11;
always @(posedge hdmi_in0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_we)
		storage_13[hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_dat_w;
	memadr_10 <= hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_11 <= hdmi2usbsoc_hdmi_in0_frame_fifo_rdport_adr;
end

assign hdmi2usbsoc_hdmi_in0_frame_fifo_wrport_dat_r = storage_13[memadr_10];
assign hdmi2usbsoc_hdmi_in0_frame_fifo_rdport_dat_r = storage_13[memadr_11];

reg [65:0] storage_14[0:15];
reg [65:0] memdat_10;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_we)
		storage_14[hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_dat_w;
	memdat_10 <= storage_14[hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_hdmi_in0_dma_fifo_wrport_dat_r = memdat_10;
assign hdmi2usbsoc_hdmi_in0_dma_fifo_rdport_dat_r = storage_14[hdmi2usbsoc_hdmi_in0_dma_fifo_rdport_adr];

reg [7:0] edid_mem_1[0:127];
reg [6:0] memadr_12;
reg [6:0] memadr_13;
always @(posedge sys_clk) begin
	memadr_12 <= hdmi2usbsoc_hdmi_in1_edid_adr;
end

always @(posedge sys_clk) begin
	if (hdmi2usbsoc_sram1_we)
		edid_mem_1[hdmi2usbsoc_sram1_adr] <= hdmi2usbsoc_sram1_dat_w;
	memadr_13 <= hdmi2usbsoc_sram1_adr;
end

assign hdmi2usbsoc_hdmi_in1_edid_dat_r = edid_mem_1[memadr_12];
assign hdmi2usbsoc_sram1_dat_r = edid_mem_1[memadr_13];

initial begin
	$readmemh("edid_mem_1.init", edid_mem_1);
end

assign hdmi_in1_sda = hdmi2usbsoc_hdmi_in1_edid_sda_drv_reg ? 1'd0 : 1'bz;
assign hdmi2usbsoc_hdmi_in1_edid_sda_i_async = hdmi_in1_sda;

IBUFDS hdmi_in_ibufds_1(
	.I(hdmi_in1_clk_p),
	.IB(hdmi_in1_clk_n),
	.O(hdmi2usbsoc_hdmi_in1_clk_input)
);

PLL_ADV #(
	.CLKFBOUT_MULT(4'd10),
	.CLKOUT0_DIVIDE(1'd1),
	.CLKOUT1_DIVIDE(3'd5),
	.CLKOUT2_DIVIDE(4'd10),
	.COMPENSATION("INTERNAL")
) hdmi_in_pll_adv_1 (
	.CLKFBIN(hdmi2usbsoc_hdmi_in1_clkfbout),
	.CLKIN1(hdmi2usbsoc_hdmi_in1_clk_input),
	.CLKINSEL(1'd1),
	.DADDR(hdmi2usbsoc_hdmi_in1_pll_adr_storage),
	.DCLK(sys_clk),
	.DEN((hdmi2usbsoc_hdmi_in1_pll_read_re | hdmi2usbsoc_hdmi_in1_pll_write_re)),
	.DI(hdmi2usbsoc_hdmi_in1_pll_dat_w_storage),
	.DWE(hdmi2usbsoc_hdmi_in1_pll_write_re),
	.RST(hdmi2usbsoc_hdmi_in1_pll_reset_storage),
	.CLKFBOUT(hdmi2usbsoc_hdmi_in1_clkfbout),
	.CLKOUT0(hdmi2usbsoc_hdmi_in1_pll_clk0),
	.CLKOUT1(hdmi2usbsoc_hdmi_in1_pll_clk1),
	.CLKOUT2(hdmi2usbsoc_hdmi_in1_pll_clk2),
	.DO(hdmi2usbsoc_hdmi_in1_pll_dat_r_status),
	.DRDY(hdmi2usbsoc_hdmi_in1_pll_drdy),
	.LOCKED(hdmi2usbsoc_hdmi_in1_pll_locked)
);

BUFPLL #(
	.DIVIDE(3'd5)
) hdmi_in_bufpll_1 (
	.GCLK(hdmi_in1_pix2x_clk),
	.LOCKED(hdmi2usbsoc_hdmi_in1_pll_locked),
	.PLLIN(hdmi2usbsoc_hdmi_in1_pll_clk0),
	.IOCLK(hdmi_in1_pix10x_clk),
	.LOCK(hdmi2usbsoc_hdmi_in1_locked_async),
	.SERDESSTROBE(hdmi2usbsoc_hdmi_in1_serdesstrobe)
);

BUFG hdmi_in_pix2x_bufg_1(
	.I(hdmi2usbsoc_hdmi_in1_pll_clk1),
	.O(hdmi_in1_pix2x_clk)
);

BUFG hdmi_in_pix_bufg_1(
	.I(hdmi2usbsoc_hdmi_in1_pll_clk2),
	.O(hdmi_in1_pix_clk)
);

IBUFDS IBUFDS_3(
	.I(hdmi_in1_data0_p),
	.IB(hdmi_in1_data0_n),
	.O(hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_se)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("STAY_AT_LIMIT"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("MASTER")
) IODELAY2_6 (
	.CAL(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_cal),
	.CE(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_ce),
	.CLK(hdmi_in1_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_se),
	.INC(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_inc),
	.IOCLK0(hdmi_in1_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_master_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_delayed_master)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("WRAPAROUND"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("SLAVE")
) IODELAY2_7 (
	.CAL(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_cal),
	.CE(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_ce),
	.CLK(hdmi_in1_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_se),
	.INC(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_inc),
	.IOCLK0(hdmi_in1_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in1_s6datacapture0_delay_slave_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_delayed_slave)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("MASTER")
) ISERDES2_22 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in1_pix10x_clk),
	.CLKDIV(hdmi_in1_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_delayed_master),
	.IOCE(hdmi2usbsoc_hdmi_in1_s6datacapture0_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_edge),
	.INCDEC(hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_incdec),
	.Q1(hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr2[1]),
	.Q2(hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr2[2]),
	.Q3(hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr2[3]),
	.Q4(hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr2[4]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_cascade),
	.VALID(hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_valid)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("SLAVE")
) ISERDES2_23 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in1_pix10x_clk),
	.CLKDIV(hdmi_in1_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in1_s6datacapture0_pad_delayed_slave),
	.IOCE(hdmi2usbsoc_hdmi_in1_s6datacapture0_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_cascade),
	.Q4(hdmi2usbsoc_hdmi_in1_s6datacapture0_dsr2[0]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in1_s6datacapture0_pd_edge)
);

IBUFDS IBUFDS_4(
	.I(hdmi_in1_data1_p),
	.IB(hdmi_in1_data1_n),
	.O(hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_se)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("STAY_AT_LIMIT"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("MASTER")
) IODELAY2_8 (
	.CAL(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_cal),
	.CE(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_ce),
	.CLK(hdmi_in1_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_se),
	.INC(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_inc),
	.IOCLK0(hdmi_in1_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_master_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_delayed_master)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("WRAPAROUND"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("SLAVE")
) IODELAY2_9 (
	.CAL(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_cal),
	.CE(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_ce),
	.CLK(hdmi_in1_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_se),
	.INC(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_inc),
	.IOCLK0(hdmi_in1_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in1_s6datacapture1_delay_slave_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_delayed_slave)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("MASTER")
) ISERDES2_24 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in1_pix10x_clk),
	.CLKDIV(hdmi_in1_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_delayed_master),
	.IOCE(hdmi2usbsoc_hdmi_in1_s6datacapture1_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_edge),
	.INCDEC(hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_incdec),
	.Q1(hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr2[1]),
	.Q2(hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr2[2]),
	.Q3(hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr2[3]),
	.Q4(hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr2[4]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_cascade),
	.VALID(hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_valid)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("SLAVE")
) ISERDES2_25 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in1_pix10x_clk),
	.CLKDIV(hdmi_in1_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in1_s6datacapture1_pad_delayed_slave),
	.IOCE(hdmi2usbsoc_hdmi_in1_s6datacapture1_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_cascade),
	.Q4(hdmi2usbsoc_hdmi_in1_s6datacapture1_dsr2[0]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in1_s6datacapture1_pd_edge)
);

IBUFDS IBUFDS_5(
	.I(hdmi_in1_data2_p),
	.IB(hdmi_in1_data2_n),
	.O(hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_se)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("STAY_AT_LIMIT"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("MASTER")
) IODELAY2_10 (
	.CAL(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_cal),
	.CE(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_ce),
	.CLK(hdmi_in1_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_se),
	.INC(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_inc),
	.IOCLK0(hdmi_in1_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_master_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_delayed_master)
);

IODELAY2 #(
	.COUNTER_WRAPAROUND("WRAPAROUND"),
	.DATA_RATE("SDR"),
	.DELAY_SRC("IDATAIN"),
	.IDELAY_TYPE("DIFF_PHASE_DETECTOR"),
	.SERDES_MODE("SLAVE")
) IODELAY2_11 (
	.CAL(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_cal),
	.CE(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_ce),
	.CLK(hdmi_in1_pix2x_clk),
	.IDATAIN(hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_se),
	.INC(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_inc),
	.IOCLK0(hdmi_in1_pix10x_clk),
	.RST(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_rst),
	.T(1'd1),
	.BUSY(hdmi2usbsoc_hdmi_in1_s6datacapture2_delay_slave_busy),
	.DATAOUT(hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_delayed_slave)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("MASTER")
) ISERDES2_26 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in1_pix10x_clk),
	.CLKDIV(hdmi_in1_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_delayed_master),
	.IOCE(hdmi2usbsoc_hdmi_in1_s6datacapture2_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_edge),
	.INCDEC(hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_incdec),
	.Q1(hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr2[1]),
	.Q2(hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr2[2]),
	.Q3(hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr2[3]),
	.Q4(hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr2[4]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_cascade),
	.VALID(hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_valid)
);

ISERDES2 #(
	.BITSLIP_ENABLE("FALSE"),
	.DATA_RATE("SDR"),
	.DATA_WIDTH(3'd5),
	.INTERFACE_TYPE("RETIMED"),
	.SERDES_MODE("SLAVE")
) ISERDES2_27 (
	.BITSLIP(1'd0),
	.CE0(1'd1),
	.CLK0(hdmi_in1_pix10x_clk),
	.CLKDIV(hdmi_in1_pix2x_clk),
	.D(hdmi2usbsoc_hdmi_in1_s6datacapture2_pad_delayed_slave),
	.IOCE(hdmi2usbsoc_hdmi_in1_s6datacapture2_serdesstrobe),
	.RST(1'd0),
	.SHIFTIN(hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_cascade),
	.Q4(hdmi2usbsoc_hdmi_in1_s6datacapture2_dsr2[0]),
	.SHIFTOUT(hdmi2usbsoc_hdmi_in1_s6datacapture2_pd_edge)
);

reg [20:0] storage_15[0:7];
reg [2:0] memadr_14;
always @(posedge hdmi_in1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_we)
		storage_15[hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_adr] <= hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_w;
	memadr_14 <= hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_adr;
end

always @(posedge hdmi_in1_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_wrport_dat_r = storage_15[memadr_14];
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_rdport_dat_r = storage_15[hdmi2usbsoc_hdmi_in1_chansync_syncbuffer0_rdport_adr];

reg [20:0] storage_16[0:7];
reg [2:0] memadr_15;
always @(posedge hdmi_in1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_we)
		storage_16[hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_adr] <= hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_w;
	memadr_15 <= hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_adr;
end

always @(posedge hdmi_in1_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_wrport_dat_r = storage_16[memadr_15];
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_rdport_dat_r = storage_16[hdmi2usbsoc_hdmi_in1_chansync_syncbuffer1_rdport_adr];

reg [20:0] storage_17[0:7];
reg [2:0] memadr_16;
always @(posedge hdmi_in1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_we)
		storage_17[hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_adr] <= hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_w;
	memadr_16 <= hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_adr;
end

always @(posedge hdmi_in1_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_wrport_dat_r = storage_17[memadr_16];
assign hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_rdport_dat_r = storage_17[hdmi2usbsoc_hdmi_in1_chansync_syncbuffer2_rdport_adr];

reg [66:0] storage_18[0:511];
reg [8:0] memadr_17;
reg [8:0] memadr_18;
always @(posedge hdmi_in1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_we)
		storage_18[hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_dat_w;
	memadr_17 <= hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_18 <= hdmi2usbsoc_hdmi_in1_frame_fifo_rdport_adr;
end

assign hdmi2usbsoc_hdmi_in1_frame_fifo_wrport_dat_r = storage_18[memadr_17];
assign hdmi2usbsoc_hdmi_in1_frame_fifo_rdport_dat_r = storage_18[memadr_18];

reg [65:0] storage_19[0:15];
reg [65:0] memdat_11;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_we)
		storage_19[hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_dat_w;
	memdat_11 <= storage_19[hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign hdmi2usbsoc_hdmi_in1_dma_fifo_wrport_dat_r = memdat_11;
assign hdmi2usbsoc_hdmi_in1_dma_fifo_rdport_dat_r = storage_19[hdmi2usbsoc_hdmi_in1_dma_fifo_rdport_adr];

reg [26:0] storage_20[0:3];
reg [1:0] memadr_19;
reg [1:0] memadr_20;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_we)
		storage_20[hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_adr] <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_dat_w;
	memadr_19 <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_20 <= hdmi2usbsoc_litedramportcdc0_cmd_fifo_rdport_adr;
end

assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_wrport_dat_r = storage_20[memadr_19];
assign hdmi2usbsoc_litedramportcdc0_cmd_fifo_rdport_dat_r = storage_20[memadr_20];

reg [65:0] storage_21[0:15];
reg [3:0] memadr_21;
reg [3:0] memadr_22;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_we)
		storage_21[hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_adr] <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_dat_w;
	memadr_21 <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	memadr_22 <= hdmi2usbsoc_litedramportcdc0_rdata_fifo_rdport_adr;
end

assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_wrport_dat_r = storage_21[memadr_21];
assign hdmi2usbsoc_litedramportcdc0_rdata_fifo_rdport_dat_r = storage_21[memadr_22];

reg [5:0] storage_22[0:3];
reg [5:0] memdat_12;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_we)
		storage_22[hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_adr] <= hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_dat_w;
	memdat_12 <= storage_22[hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_adr];
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_wrport_dat_r = memdat_12;
assign hdmi2usbsoc_litedramportconverter0_cmd_buffer_rdport_dat_r = storage_22[hdmi2usbsoc_litedramportconverter0_cmd_buffer_rdport_adr];

reg [161:0] storage_23[0:1];
reg [0:0] memadr_23;
reg [0:0] memadr_24;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_we)
		storage_23[hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_adr] <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_dat_w;
	memadr_23 <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	memadr_24 <= hdmi2usbsoc_hdmi_out0_core_initiator_cdc_rdport_adr;
end

assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_wrport_dat_r = storage_23[memadr_23];
assign hdmi2usbsoc_hdmi_out0_core_initiator_cdc_rdport_dat_r = storage_23[memadr_24];

reg [17:0] storage_24[0:4095];
reg [17:0] memdat_13;
reg [17:0] memdat_14;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_we)
		storage_24[hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_dat_w;
	memdat_13 <= storage_24[hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_adr];
end

always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_re)
		memdat_14 <= storage_24[hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_adr];
end

assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_wrport_dat_r = memdat_13;
assign hdmi2usbsoc_hdmi_out0_core_dmareader_fifo_rdport_dat_r = memdat_14;

DCM_CLKGEN #(
	.CLKFXDV_DIVIDE(2'd2),
	.CLKFX_DIVIDE(3'd4),
	.CLKFX_MD_MAX(2.0),
	.CLKFX_MULTIPLY(2'd2),
	.CLKIN_PERIOD(20.0),
	.SPREAD_SPECTRUM("NONE"),
	.STARTUP_WAIT("FALSE")
) hdmi_out_dcm_clkgen (
	.CLKIN(base50_clk),
	.FREEZEDCM(1'd0),
	.PROGCLK(sys_clk),
	.PROGDATA(hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progdata),
	.PROGEN(hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progen),
	.RST(sys_rst),
	.CLKFX(hdmi2usbsoc_hdmi_out0_driver_clocking_clk_pix_unbuffered),
	.LOCKED(hdmi2usbsoc_hdmi_out0_driver_clocking_pix_locked),
	.PROGDONE(hdmi2usbsoc_hdmi_out0_driver_clocking_pix_progdone)
);

PLL_ADV #(
	.CLKFBOUT_MULT(4'd10),
	.CLKOUT0_DIVIDE(1'd1),
	.CLKOUT1_DIVIDE(3'd5),
	.CLKOUT2_DIVIDE(4'd10),
	.COMPENSATION("INTERNAL")
) hdmi_out_pll_adv (
	.CLKFBIN(hdmi2usbsoc_hdmi_out0_driver_clocking_clkfbout),
	.CLKIN1(hdmi2usbsoc_hdmi_out0_driver_clocking_clk_pix_unbuffered),
	.CLKINSEL(1'd1),
	.DADDR(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_adr_storage),
	.DCLK(sys_clk),
	.DEN((hdmi2usbsoc_hdmi_out0_driver_clocking_pll_read_re | hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_re)),
	.DI(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_w_storage),
	.DWE(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_write_re),
	.RST(((~hdmi2usbsoc_hdmi_out0_driver_clocking_pix_locked) | hdmi2usbsoc_hdmi_out0_driver_clocking_pll_reset_storage)),
	.CLKFBOUT(hdmi2usbsoc_hdmi_out0_driver_clocking_clkfbout),
	.CLKOUT0(hdmi2usbsoc_hdmi_out0_driver_clocking_pll0_pix10x),
	.CLKOUT1(hdmi2usbsoc_hdmi_out0_driver_clocking_pll1_pix2x),
	.CLKOUT2(hdmi2usbsoc_hdmi_out0_driver_clocking_pll2_pix),
	.DO(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_dat_r_status),
	.DRDY(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_drdy),
	.LOCKED(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_locked)
);

BUFPLL #(
	.DIVIDE(3'd5)
) hdmi_out_bufpll (
	.GCLK(hdmi_out0_pix2x_clk),
	.LOCKED(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_locked),
	.PLLIN(hdmi2usbsoc_hdmi_out0_driver_clocking_pll0_pix10x),
	.IOCLK(hdmi_out0_pix10x_clk),
	.LOCK(hdmi2usbsoc_hdmi_out0_driver_clocking_locked_async),
	.SERDESSTROBE(hdmi2usbsoc_hdmi_out0_driver_clocking_serdesstrobe)
);

BUFG hdmi_out_pix2x_bufg(
	.I(hdmi2usbsoc_hdmi_out0_driver_clocking_pll1_pix2x),
	.O(hdmi_out0_pix2x_clk)
);

BUFG hdmi_out_pix_bufg(
	.I(hdmi2usbsoc_hdmi_out0_driver_clocking_pll2_pix),
	.O(hdmi_out0_pix_clk)
);

ODDR2 #(
	.DDR_ALIGNMENT("NONE"),
	.INIT(1'd0),
	.SRTYPE("SYNC")
) ODDR2_5 (
	.C0(hdmi_out0_pix_clk),
	.C1((~hdmi_out0_pix_clk)),
	.CE(1'd1),
	.D0(1'd1),
	.D1(1'd0),
	.R(1'd0),
	.S(1'd0),
	.Q(hdmi2usbsoc_hdmi_out0_driver_clocking_hdmi_clk_se)
);

OBUFDS OBUFDS_1(
	.I(hdmi2usbsoc_hdmi_out0_driver_clocking_hdmi_clk_se),
	.O(hdmi_out0_clk_p),
	.OB(hdmi_out0_clk_n)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("MASTER")
) OSERDES2_18 (
	.CLK0(hdmi_out0_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out0_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x[4]),
	.D2(1'd0),
	.D3(1'd0),
	.D4(1'd0),
	.IOCE(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd1),
	.SHIFTIN2(1'd1),
	.SHIFTIN3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_do),
	.SHIFTIN4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_to),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_pad_se),
	.SHIFTOUT1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_di),
	.SHIFTOUT2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_ti)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("SLAVE")
) OSERDES2_19 (
	.CLK0(hdmi_out0_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out0_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x[0]),
	.D2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x[1]),
	.D3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x[2]),
	.D4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_ed_2x[3]),
	.IOCE(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_di),
	.SHIFTIN2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_ti),
	.SHIFTIN3(1'd1),
	.SHIFTIN4(1'd1),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.SHIFTOUT3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_do),
	.SHIFTOUT4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_cascade_to)
);

OBUFDS OBUFDS_2(
	.I(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es0_pad_se),
	.O(hdmi_out0_data0_p),
	.OB(hdmi_out0_data0_n)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("MASTER")
) OSERDES2_20 (
	.CLK0(hdmi_out0_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out0_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x[4]),
	.D2(1'd0),
	.D3(1'd0),
	.D4(1'd0),
	.IOCE(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd1),
	.SHIFTIN2(1'd1),
	.SHIFTIN3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_do),
	.SHIFTIN4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_to),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_pad_se),
	.SHIFTOUT1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_di),
	.SHIFTOUT2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_ti)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("SLAVE")
) OSERDES2_21 (
	.CLK0(hdmi_out0_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out0_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x[0]),
	.D2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x[1]),
	.D3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x[2]),
	.D4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_ed_2x[3]),
	.IOCE(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_di),
	.SHIFTIN2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_ti),
	.SHIFTIN3(1'd1),
	.SHIFTIN4(1'd1),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.SHIFTOUT3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_do),
	.SHIFTOUT4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_cascade_to)
);

OBUFDS OBUFDS_3(
	.I(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es1_pad_se),
	.O(hdmi_out0_data1_p),
	.OB(hdmi_out0_data1_n)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("MASTER")
) OSERDES2_22 (
	.CLK0(hdmi_out0_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out0_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x[4]),
	.D2(1'd0),
	.D3(1'd0),
	.D4(1'd0),
	.IOCE(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd1),
	.SHIFTIN2(1'd1),
	.SHIFTIN3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_do),
	.SHIFTIN4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_to),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_pad_se),
	.SHIFTOUT1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_di),
	.SHIFTOUT2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_ti)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("SLAVE")
) OSERDES2_23 (
	.CLK0(hdmi_out0_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out0_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x[0]),
	.D2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x[1]),
	.D3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x[2]),
	.D4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_ed_2x[3]),
	.IOCE(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_di),
	.SHIFTIN2(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_ti),
	.SHIFTIN3(1'd1),
	.SHIFTIN4(1'd1),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.SHIFTOUT3(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_do),
	.SHIFTOUT4(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_cascade_to)
);

OBUFDS OBUFDS_4(
	.I(hdmi2usbsoc_hdmi_out0_driver_hdmi_phy_es2_pad_se),
	.O(hdmi_out0_data2_p),
	.OB(hdmi_out0_data2_n)
);

reg [9:0] storage_25[0:3];
reg [9:0] memdat_15;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_we)
		storage_25[hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_dat_w;
	memdat_15 <= storage_25[hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_adr];
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_wrport_dat_r = memdat_15;
assign hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_rdport_dat_r = storage_25[hdmi2usbsoc_hdmi_out0_resetinserter_y_fifo_rdport_adr];

reg [9:0] storage_26[0:3];
reg [9:0] memdat_16;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_we)
		storage_26[hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_w;
	memdat_16 <= storage_26[hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_adr];
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_r = memdat_16;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_rdport_dat_r = storage_26[hdmi2usbsoc_hdmi_out0_resetinserter_cb_fifo_rdport_adr];

reg [9:0] storage_27[0:3];
reg [9:0] memdat_17;
always @(posedge hdmi_out0_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_we)
		storage_27[hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_w;
	memdat_17 <= storage_27[hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_adr];
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_r = memdat_17;
assign hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_rdport_dat_r = storage_27[hdmi2usbsoc_hdmi_out0_resetinserter_cr_fifo_rdport_adr];

reg [26:0] storage_28[0:3];
reg [1:0] memadr_25;
reg [1:0] memadr_26;
always @(posedge hdmi_out1_pix_clk) begin
	if (hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_we)
		storage_28[hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_adr] <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_dat_w;
	memadr_25 <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_26 <= hdmi2usbsoc_litedramportcdc1_cmd_fifo_rdport_adr;
end

assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_wrport_dat_r = storage_28[memadr_25];
assign hdmi2usbsoc_litedramportcdc1_cmd_fifo_rdport_dat_r = storage_28[memadr_26];

reg [65:0] storage_29[0:15];
reg [3:0] memadr_27;
reg [3:0] memadr_28;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_we)
		storage_29[hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_adr] <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_dat_w;
	memadr_27 <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_adr;
end

always @(posedge hdmi_out1_pix_clk) begin
	memadr_28 <= hdmi2usbsoc_litedramportcdc1_rdata_fifo_rdport_adr;
end

assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_wrport_dat_r = storage_29[memadr_27];
assign hdmi2usbsoc_litedramportcdc1_rdata_fifo_rdport_dat_r = storage_29[memadr_28];

reg [5:0] storage_30[0:3];
reg [5:0] memdat_18;
always @(posedge hdmi_out1_pix_clk) begin
	if (hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_we)
		storage_30[hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_adr] <= hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_dat_w;
	memdat_18 <= storage_30[hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_adr];
end

always @(posedge hdmi_out1_pix_clk) begin
end

assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_wrport_dat_r = memdat_18;
assign hdmi2usbsoc_litedramportconverter1_cmd_buffer_rdport_dat_r = storage_30[hdmi2usbsoc_litedramportconverter1_cmd_buffer_rdport_adr];

reg [161:0] storage_31[0:1];
reg [0:0] memadr_29;
reg [0:0] memadr_30;
always @(posedge sys_clk) begin
	if (hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_we)
		storage_31[hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_adr] <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_dat_w;
	memadr_29 <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_adr;
end

always @(posedge hdmi_out1_pix_clk) begin
	memadr_30 <= hdmi2usbsoc_hdmi_out1_core_initiator_cdc_rdport_adr;
end

assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_wrport_dat_r = storage_31[memadr_29];
assign hdmi2usbsoc_hdmi_out1_core_initiator_cdc_rdport_dat_r = storage_31[memadr_30];

reg [17:0] storage_32[0:4095];
reg [17:0] memdat_19;
reg [17:0] memdat_20;
always @(posedge hdmi_out1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_we)
		storage_32[hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_dat_w;
	memdat_19 <= storage_32[hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_adr];
end

always @(posedge hdmi_out1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_re)
		memdat_20 <= storage_32[hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_adr];
end

assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_wrport_dat_r = memdat_19;
assign hdmi2usbsoc_hdmi_out1_core_dmareader_fifo_rdport_dat_r = memdat_20;

BUFG hdmi_out_pix_bufg_1(
	.I(hdmi2usbsoc_hdmi_out0_driver_clocking_pll2_pix),
	.O(hdmi_out1_pix_clk)
);

BUFG hdmi_out_pix2x_bufg_1(
	.I(hdmi2usbsoc_hdmi_out0_driver_clocking_pll1_pix2x),
	.O(hdmi_out1_pix2x_clk)
);

BUFPLL #(
	.DIVIDE(3'd5)
) hdmi_out_bufpll_1 (
	.GCLK(hdmi_out1_pix2x_clk),
	.LOCKED(hdmi2usbsoc_hdmi_out0_driver_clocking_pll_locked),
	.PLLIN(hdmi2usbsoc_hdmi_out0_driver_clocking_pll0_pix10x),
	.IOCLK(hdmi_out1_pix10x_clk),
	.SERDESSTROBE(hdmi2usbsoc_hdmi_out1_driver_clocking_serdesstrobe)
);

ODDR2 #(
	.DDR_ALIGNMENT("NONE"),
	.INIT(1'd0),
	.SRTYPE("SYNC")
) ODDR2_6 (
	.C0(hdmi_out1_pix_clk),
	.C1((~hdmi_out1_pix_clk)),
	.CE(1'd1),
	.D0(1'd1),
	.D1(1'd0),
	.R(1'd0),
	.S(1'd0),
	.Q(hdmi2usbsoc_hdmi_out1_driver_clocking_hdmi_clk_se)
);

OBUFDS OBUFDS_5(
	.I(hdmi2usbsoc_hdmi_out1_driver_clocking_hdmi_clk_se),
	.O(hdmi_out1_clk_p),
	.OB(hdmi_out1_clk_n)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("MASTER")
) OSERDES2_24 (
	.CLK0(hdmi_out1_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out1_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x[4]),
	.D2(1'd0),
	.D3(1'd0),
	.D4(1'd0),
	.IOCE(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd1),
	.SHIFTIN2(1'd1),
	.SHIFTIN3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_do),
	.SHIFTIN4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_to),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_pad_se),
	.SHIFTOUT1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_di),
	.SHIFTOUT2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_ti)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("SLAVE")
) OSERDES2_25 (
	.CLK0(hdmi_out1_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out1_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x[0]),
	.D2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x[1]),
	.D3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x[2]),
	.D4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_ed_2x[3]),
	.IOCE(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_di),
	.SHIFTIN2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_ti),
	.SHIFTIN3(1'd1),
	.SHIFTIN4(1'd1),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.SHIFTOUT3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_do),
	.SHIFTOUT4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_cascade_to)
);

OBUFDS OBUFDS_6(
	.I(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es0_pad_se),
	.O(hdmi_out1_data0_p),
	.OB(hdmi_out1_data0_n)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("MASTER")
) OSERDES2_26 (
	.CLK0(hdmi_out1_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out1_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x[4]),
	.D2(1'd0),
	.D3(1'd0),
	.D4(1'd0),
	.IOCE(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd1),
	.SHIFTIN2(1'd1),
	.SHIFTIN3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_do),
	.SHIFTIN4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_to),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_pad_se),
	.SHIFTOUT1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_di),
	.SHIFTOUT2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_ti)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("SLAVE")
) OSERDES2_27 (
	.CLK0(hdmi_out1_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out1_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x[0]),
	.D2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x[1]),
	.D3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x[2]),
	.D4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_ed_2x[3]),
	.IOCE(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_di),
	.SHIFTIN2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_ti),
	.SHIFTIN3(1'd1),
	.SHIFTIN4(1'd1),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.SHIFTOUT3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_do),
	.SHIFTOUT4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_cascade_to)
);

OBUFDS OBUFDS_7(
	.I(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es1_pad_se),
	.O(hdmi_out1_data1_p),
	.OB(hdmi_out1_data1_n)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("MASTER")
) OSERDES2_28 (
	.CLK0(hdmi_out1_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out1_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x[4]),
	.D2(1'd0),
	.D3(1'd0),
	.D4(1'd0),
	.IOCE(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(1'd1),
	.SHIFTIN2(1'd1),
	.SHIFTIN3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_do),
	.SHIFTIN4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_to),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.OQ(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_pad_se),
	.SHIFTOUT1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_di),
	.SHIFTOUT2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_ti)
);

OSERDES2 #(
	.DATA_RATE_OQ("SDR"),
	.DATA_RATE_OT("SDR"),
	.DATA_WIDTH(3'd5),
	.OUTPUT_MODE("DIFFERENTIAL"),
	.SERDES_MODE("SLAVE")
) OSERDES2_29 (
	.CLK0(hdmi_out1_pix10x_clk),
	.CLK1(1'd0),
	.CLKDIV(hdmi_out1_pix2x_clk),
	.D1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x[0]),
	.D2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x[1]),
	.D3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x[2]),
	.D4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_ed_2x[3]),
	.IOCE(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_serdesstrobe),
	.OCE(1'd1),
	.RST(1'd0),
	.SHIFTIN1(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_di),
	.SHIFTIN2(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_ti),
	.SHIFTIN3(1'd1),
	.SHIFTIN4(1'd1),
	.T1(1'd0),
	.T2(1'd0),
	.T3(1'd0),
	.T4(1'd0),
	.TCE(1'd1),
	.TRAIN(1'd0),
	.SHIFTOUT3(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_do),
	.SHIFTOUT4(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_cascade_to)
);

OBUFDS OBUFDS_8(
	.I(hdmi2usbsoc_hdmi_out1_driver_hdmi_phy_es2_pad_se),
	.O(hdmi_out1_data2_p),
	.OB(hdmi_out1_data2_n)
);

reg [9:0] storage_33[0:3];
reg [9:0] memdat_21;
always @(posedge hdmi_out1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_we)
		storage_33[hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_dat_w;
	memdat_21 <= storage_33[hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_adr];
end

always @(posedge hdmi_out1_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_wrport_dat_r = memdat_21;
assign hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_rdport_dat_r = storage_33[hdmi2usbsoc_hdmi_out1_resetinserter_y_fifo_rdport_adr];

reg [9:0] storage_34[0:3];
reg [9:0] memdat_22;
always @(posedge hdmi_out1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_we)
		storage_34[hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_dat_w;
	memdat_22 <= storage_34[hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_adr];
end

always @(posedge hdmi_out1_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_wrport_dat_r = memdat_22;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_rdport_dat_r = storage_34[hdmi2usbsoc_hdmi_out1_resetinserter_cb_fifo_rdport_adr];

reg [9:0] storage_35[0:3];
reg [9:0] memdat_23;
always @(posedge hdmi_out1_pix_clk) begin
	if (hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_we)
		storage_35[hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_adr] <= hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_dat_w;
	memdat_23 <= storage_35[hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_adr];
end

always @(posedge hdmi_out1_pix_clk) begin
end

assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_wrport_dat_r = memdat_23;
assign hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_rdport_dat_r = storage_35[hdmi2usbsoc_hdmi_out1_resetinserter_cr_fifo_rdport_adr];

reg [129:0] storage_36[0:15];
reg [129:0] memdat_24;
always @(posedge sys_clk) begin
	if (encoder_reader_fifo_wrport_we)
		storage_36[encoder_reader_fifo_wrport_adr] <= encoder_reader_fifo_wrport_dat_w;
	memdat_24 <= storage_36[encoder_reader_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign encoder_reader_fifo_wrport_dat_r = memdat_24;
assign encoder_reader_fifo_rdport_dat_r = storage_36[encoder_reader_fifo_rdport_adr];

reg [129:0] storage_37[0:3];
reg [1:0] memadr_31;
reg [1:0] memadr_32;
always @(posedge sys_clk) begin
	if (encoder_cdc_wrport_we)
		storage_37[encoder_cdc_wrport_adr] <= encoder_cdc_wrport_dat_w;
	memadr_31 <= encoder_cdc_wrport_adr;
end

always @(posedge encoder_clk) begin
	memadr_32 <= encoder_cdc_rdport_adr;
end

assign encoder_cdc_wrport_dat_r = storage_37[memadr_31];
assign encoder_cdc_rdport_dat_r = storage_37[memadr_32];

reg [127:0] mem_3[0:15];
reg [3:0] memadr_33;
always @(posedge encoder_clk) begin
	if (encoderbuffer_write_port_we)
		mem_3[encoderbuffer_write_port_adr] <= encoderbuffer_write_port_dat_w;
	memadr_33 <= encoderbuffer_write_port_adr;
end

always @(posedge encoder_clk) begin
end

assign encoderbuffer_write_port_dat_r = mem_3[memadr_33];
assign encoderbuffer_read_port_dat_r = mem_3[encoderbuffer_read_port_adr];

reg [9:0] storage_38[0:3];
reg [9:0] memdat_25;
always @(posedge encoder_clk) begin
	if (encoder_y_fifo_wrport_we)
		storage_38[encoder_y_fifo_wrport_adr] <= encoder_y_fifo_wrport_dat_w;
	memdat_25 <= storage_38[encoder_y_fifo_wrport_adr];
end

always @(posedge encoder_clk) begin
end

assign encoder_y_fifo_wrport_dat_r = memdat_25;
assign encoder_y_fifo_rdport_dat_r = storage_38[encoder_y_fifo_rdport_adr];

reg [9:0] storage_39[0:3];
reg [9:0] memdat_26;
always @(posedge encoder_clk) begin
	if (encoder_cb_fifo_wrport_we)
		storage_39[encoder_cb_fifo_wrport_adr] <= encoder_cb_fifo_wrport_dat_w;
	memdat_26 <= storage_39[encoder_cb_fifo_wrport_adr];
end

always @(posedge encoder_clk) begin
end

assign encoder_cb_fifo_wrport_dat_r = memdat_26;
assign encoder_cb_fifo_rdport_dat_r = storage_39[encoder_cb_fifo_rdport_adr];

reg [9:0] storage_40[0:3];
reg [9:0] memdat_27;
always @(posedge encoder_clk) begin
	if (encoder_cr_fifo_wrport_we)
		storage_40[encoder_cr_fifo_wrport_adr] <= encoder_cr_fifo_wrport_dat_w;
	memdat_27 <= storage_40[encoder_cr_fifo_wrport_adr];
end

always @(posedge encoder_clk) begin
end

assign encoder_cr_fifo_wrport_dat_r = memdat_27;
assign encoder_cr_fifo_rdport_dat_r = storage_40[encoder_cr_fifo_rdport_adr];

reg [9:0] storage_41[0:1023];
reg [9:0] memdat_28;
reg [9:0] memdat_29;
always @(posedge encoder_clk) begin
	if (encoder_output_fifo_wrport_we)
		storage_41[encoder_output_fifo_wrport_adr] <= encoder_output_fifo_wrport_dat_w;
	memdat_28 <= storage_41[encoder_output_fifo_wrport_adr];
end

always @(posedge encoder_clk) begin
	if (encoder_output_fifo_rdport_re)
		memdat_29 <= storage_41[encoder_output_fifo_rdport_adr];
end

assign encoder_output_fifo_wrport_dat_r = memdat_28;
assign encoder_output_fifo_rdport_dat_r = memdat_29;

wb_async_reg wb_async_reg(
	.wbm_adr_i(encoder_bus_adr),
	.wbm_clk(sys_clk),
	.wbm_cyc_i(encoder_bus_cyc),
	.wbm_dat_i(encoder_bus_dat_w),
	.wbm_rst(sys_rst),
	.wbm_sel_i(encoder_bus_sel),
	.wbm_stb_i(encoder_bus_stb),
	.wbm_we_i(encoder_bus_we),
	.wbs_ack_i(encoder_jpeg_bus_ack),
	.wbs_clk(encoder_clk),
	.wbs_dat_i(encoder_jpeg_bus_dat_r),
	.wbs_err_i(encoder_jpeg_bus_err),
	.wbs_rst(encoder_rst),
	.wbs_rty_i(1'd0),
	.wbm_ack_o(encoder_bus_ack),
	.wbm_dat_o(encoder_bus_dat_r),
	.wbm_err_o(encoder_bus_err),
	.wbs_adr_o(encoder_jpeg_bus_adr),
	.wbs_cyc_o(encoder_jpeg_bus_cyc),
	.wbs_dat_o(encoder_jpeg_bus_dat_w),
	.wbs_sel_o(encoder_jpeg_bus_sel),
	.wbs_stb_o(encoder_jpeg_bus_stb),
	.wbs_we_o(encoder_jpeg_bus_we)
);

JpegEnc JpegEnc(
	.CLK(encoder_clk),
	.OPB_ABus(({encoder_jpeg_bus_adr, encoder} & 10'd1023)),
	.OPB_BE(encoder_jpeg_bus_sel),
	.OPB_DBus_in(encoder_jpeg_bus_dat_w),
	.OPB_RNW((~encoder_jpeg_bus_we)),
	.OPB_select((encoder_jpeg_bus_stb & encoder_jpeg_bus_cyc)),
	.RST(encoder_rst),
	.fdct_fifo_hf_full(encoder_fdct_fifo_hf_full),
	.fdct_fifo_q(encoder_fdct_fifo_q),
	.outif_almost_full(encoder_output_fifo_almost_full),
	.OPB_DBus_out(encoder_jpeg_bus_dat_r),
	.OPB_XferAck(encoder_jpeg_bus_ack),
	.OPB_errAck(encoder_jpeg_bus_err),
	.fdct_fifo_rd(encoder_fdct_fifo_rd),
	.ram_byte(encoder_output_fifo_sink_payload_data),
	.ram_wren(encoder_output_fifo_sink_valid)
);

IBUFG IBUFG_1(
	.I(fx2_ifclk),
	.O(usb_clk)
);

reg [9:0] storage_42[0:3];
reg [1:0] memadr_34;
reg [1:0] memadr_35;
always @(posedge encoder_clk) begin
	if (encoder_streamer_fifo_wrport_we)
		storage_42[encoder_streamer_fifo_wrport_adr] <= encoder_streamer_fifo_wrport_dat_w;
	memadr_34 <= encoder_streamer_fifo_wrport_adr;
end

always @(posedge usb_clk) begin
	memadr_35 <= encoder_streamer_fifo_rdport_adr;
end

assign encoder_streamer_fifo_wrport_dat_r = storage_42[memadr_34];
assign encoder_streamer_fifo_rdport_dat_r = storage_42[memadr_35];

fx2_jpeg_streamer fx2_jpeg_streamer(
	.clk(usb_clk),
	.fx2_empty_n(fx2_flagc),
	.fx2_full_n(fx2_flagb),
	.rst(usb_rst),
	.sink_data(encoder_streamer_fifo_source_payload_data),
	.sink_stb(encoder_streamer_fifo_source_valid),
	.fx2_data(fx2_data),
	.fx2_addr(fx2_addr),
	.fx2_cs_n(fx2_cs_n),
	.fx2_oe_n(fx2_oe_n),
	.fx2_pktend_n(fx2_pktend_n),
	.fx2_rd_n(fx2_rd_n),
	.fx2_wr_n(fx2_wr_n),
	.sink_ack(encoder_streamer_fifo_source_ready)
);

FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(por_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl0),
	.Q(xilinxasyncresetsynchronizerimpl0_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(por_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl0),
	.Q(por_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl1),
	.Q(xilinxasyncresetsynchronizerimpl1_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(sys_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl1),
	.Q(sys_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(base50_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl2),
	.Q(xilinxasyncresetsynchronizerimpl2_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(base50_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl2),
	.Q(base50_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(encoder_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(sys_rst),
	.Q(xilinxasyncresetsynchronizerimpl3_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(encoder_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(sys_rst),
	.Q(encoder_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_8 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl4),
	.Q(xilinxasyncresetsynchronizerimpl4_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_9 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl4_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl4),
	.Q(hdmi_in0_pix_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_10 (
	.C(hdmi_in0_pix2x_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl5),
	.Q(xilinxasyncresetsynchronizerimpl5_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_11 (
	.C(hdmi_in0_pix2x_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl5_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl5),
	.Q(hdmi_in0_pix2x_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_12 (
	.C(hdmi_in1_pix_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl6),
	.Q(xilinxasyncresetsynchronizerimpl6_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_13 (
	.C(hdmi_in1_pix_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl6_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl6),
	.Q(hdmi_in1_pix_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_14 (
	.C(hdmi_in1_pix2x_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(xilinxasyncresetsynchronizerimpl7),
	.Q(xilinxasyncresetsynchronizerimpl7_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_15 (
	.C(hdmi_in1_pix2x_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl7_rst_meta),
	.PRE(xilinxasyncresetsynchronizerimpl7),
	.Q(hdmi_in1_pix2x_rst)
);

FDPE #(
	.INIT(1'd1)
) FDPE_16 (
	.C(usb_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(sys_rst),
	.Q(xilinxasyncresetsynchronizerimpl8_rst_meta)
);

FDPE #(
	.INIT(1'd1)
) FDPE_17 (
	.C(usb_clk),
	.CE(1'd1),
	.D(xilinxasyncresetsynchronizerimpl8_rst_meta),
	.PRE(sys_rst),
	.Q(usb_rst)
);

endmodule
